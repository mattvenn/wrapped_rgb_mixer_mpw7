// This is the unpowered netlist.
module wrapped_rgb_mixer (active,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la1_data_in,
    la1_data_out,
    la1_oenb);
 input active;
 input wb_clk_i;
 input [37:0] io_in;
 inout [37:0] io_oeb;
 inout [37:0] io_out;
 input [31:0] la1_data_in;
 inout [31:0] la1_data_out;
 input [31:0] la1_oenb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire clknet_0_wb_clk_i;
 wire \rgb_mixer.debounce0_a.button_hist[0] ;
 wire \rgb_mixer.debounce0_a.button_hist[1] ;
 wire \rgb_mixer.debounce0_a.button_hist[2] ;
 wire \rgb_mixer.debounce0_a.button_hist[3] ;
 wire \rgb_mixer.debounce0_a.button_hist[4] ;
 wire \rgb_mixer.debounce0_a.button_hist[5] ;
 wire \rgb_mixer.debounce0_a.button_hist[6] ;
 wire \rgb_mixer.debounce0_a.button_hist[7] ;
 wire \rgb_mixer.debounce0_a.debounced ;
 wire \rgb_mixer.debounce0_b.button_hist[0] ;
 wire \rgb_mixer.debounce0_b.button_hist[1] ;
 wire \rgb_mixer.debounce0_b.button_hist[2] ;
 wire \rgb_mixer.debounce0_b.button_hist[3] ;
 wire \rgb_mixer.debounce0_b.button_hist[4] ;
 wire \rgb_mixer.debounce0_b.button_hist[5] ;
 wire \rgb_mixer.debounce0_b.button_hist[6] ;
 wire \rgb_mixer.debounce0_b.button_hist[7] ;
 wire \rgb_mixer.debounce0_b.debounced ;
 wire \rgb_mixer.debounce1_a.button_hist[0] ;
 wire \rgb_mixer.debounce1_a.button_hist[1] ;
 wire \rgb_mixer.debounce1_a.button_hist[2] ;
 wire \rgb_mixer.debounce1_a.button_hist[3] ;
 wire \rgb_mixer.debounce1_a.button_hist[4] ;
 wire \rgb_mixer.debounce1_a.button_hist[5] ;
 wire \rgb_mixer.debounce1_a.button_hist[6] ;
 wire \rgb_mixer.debounce1_a.button_hist[7] ;
 wire \rgb_mixer.debounce1_a.debounced ;
 wire \rgb_mixer.debounce1_b.button_hist[0] ;
 wire \rgb_mixer.debounce1_b.button_hist[1] ;
 wire \rgb_mixer.debounce1_b.button_hist[2] ;
 wire \rgb_mixer.debounce1_b.button_hist[3] ;
 wire \rgb_mixer.debounce1_b.button_hist[4] ;
 wire \rgb_mixer.debounce1_b.button_hist[5] ;
 wire \rgb_mixer.debounce1_b.button_hist[6] ;
 wire \rgb_mixer.debounce1_b.button_hist[7] ;
 wire \rgb_mixer.debounce1_b.debounced ;
 wire \rgb_mixer.debounce2_a.button_hist[0] ;
 wire \rgb_mixer.debounce2_a.button_hist[1] ;
 wire \rgb_mixer.debounce2_a.button_hist[2] ;
 wire \rgb_mixer.debounce2_a.button_hist[3] ;
 wire \rgb_mixer.debounce2_a.button_hist[4] ;
 wire \rgb_mixer.debounce2_a.button_hist[5] ;
 wire \rgb_mixer.debounce2_a.button_hist[6] ;
 wire \rgb_mixer.debounce2_a.button_hist[7] ;
 wire \rgb_mixer.debounce2_a.debounced ;
 wire \rgb_mixer.debounce2_b.button_hist[0] ;
 wire \rgb_mixer.debounce2_b.button_hist[1] ;
 wire \rgb_mixer.debounce2_b.button_hist[2] ;
 wire \rgb_mixer.debounce2_b.button_hist[3] ;
 wire \rgb_mixer.debounce2_b.button_hist[4] ;
 wire \rgb_mixer.debounce2_b.button_hist[5] ;
 wire \rgb_mixer.debounce2_b.button_hist[6] ;
 wire \rgb_mixer.debounce2_b.button_hist[7] ;
 wire \rgb_mixer.debounce2_b.debounced ;
 wire \rgb_mixer.enc0[0] ;
 wire \rgb_mixer.enc0[1] ;
 wire \rgb_mixer.enc0[2] ;
 wire \rgb_mixer.enc0[3] ;
 wire \rgb_mixer.enc0[4] ;
 wire \rgb_mixer.enc0[5] ;
 wire \rgb_mixer.enc0[6] ;
 wire \rgb_mixer.enc0[7] ;
 wire \rgb_mixer.enc1[0] ;
 wire \rgb_mixer.enc1[1] ;
 wire \rgb_mixer.enc1[2] ;
 wire \rgb_mixer.enc1[3] ;
 wire \rgb_mixer.enc1[4] ;
 wire \rgb_mixer.enc1[5] ;
 wire \rgb_mixer.enc1[6] ;
 wire \rgb_mixer.enc1[7] ;
 wire \rgb_mixer.enc2[0] ;
 wire \rgb_mixer.enc2[1] ;
 wire \rgb_mixer.enc2[2] ;
 wire \rgb_mixer.enc2[3] ;
 wire \rgb_mixer.enc2[4] ;
 wire \rgb_mixer.enc2[5] ;
 wire \rgb_mixer.enc2[6] ;
 wire \rgb_mixer.enc2[7] ;
 wire \rgb_mixer.encoder0.old_a ;
 wire \rgb_mixer.encoder0.old_b ;
 wire \rgb_mixer.encoder1.old_a ;
 wire \rgb_mixer.encoder1.old_b ;
 wire \rgb_mixer.encoder2.old_a ;
 wire \rgb_mixer.encoder2.old_b ;
 wire \rgb_mixer.pwm0.count[0] ;
 wire \rgb_mixer.pwm0.count[1] ;
 wire \rgb_mixer.pwm0.count[2] ;
 wire \rgb_mixer.pwm0.count[3] ;
 wire \rgb_mixer.pwm0.count[4] ;
 wire \rgb_mixer.pwm0.count[5] ;
 wire \rgb_mixer.pwm0.count[6] ;
 wire \rgb_mixer.pwm0.count[7] ;
 wire \rgb_mixer.pwm0.out ;
 wire \rgb_mixer.pwm1.count[0] ;
 wire \rgb_mixer.pwm1.count[1] ;
 wire \rgb_mixer.pwm1.count[2] ;
 wire \rgb_mixer.pwm1.count[3] ;
 wire \rgb_mixer.pwm1.count[4] ;
 wire \rgb_mixer.pwm1.count[5] ;
 wire \rgb_mixer.pwm1.count[6] ;
 wire \rgb_mixer.pwm1.count[7] ;
 wire \rgb_mixer.pwm1.out ;
 wire \rgb_mixer.pwm2.count[0] ;
 wire \rgb_mixer.pwm2.count[1] ;
 wire \rgb_mixer.pwm2.count[2] ;
 wire \rgb_mixer.pwm2.count[3] ;
 wire \rgb_mixer.pwm2.count[4] ;
 wire \rgb_mixer.pwm2.count[5] ;
 wire \rgb_mixer.pwm2.count[6] ;
 wire \rgb_mixer.pwm2.count[7] ;
 wire \rgb_mixer.pwm2.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 sky130_fd_sc_hd__buf_6 _0663_ (.A(net1),
    .X(_0108_));
 sky130_fd_sc_hd__buf_12 _0664_ (.A(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_8 _0665_ (.A(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__inv_2 _0666_ (.A(_0110_),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _0667_ (.A(_0110_),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _0668_ (.A(_0110_),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_2 _0669_ (.A(_0110_),
    .Y(_0460_));
 sky130_fd_sc_hd__inv_2 _0670_ (.A(_0110_),
    .Y(_0459_));
 sky130_fd_sc_hd__inv_2 _0671_ (.A(_0110_),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_2 _0672_ (.A(_0110_),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(_0110_),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(_0110_),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(_0110_),
    .Y(_0463_));
 sky130_fd_sc_hd__buf_8 _0676_ (.A(_0109_),
    .X(_0111_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(_0111_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _0678_ (.A(_0111_),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_2 _0679_ (.A(_0111_),
    .Y(_0455_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(_0111_),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _0681_ (.A(_0111_),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(_0111_),
    .Y(_0467_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(_0111_),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(_0111_),
    .Y(_0469_));
 sky130_fd_sc_hd__inv_2 _0685_ (.A(_0111_),
    .Y(_0470_));
 sky130_fd_sc_hd__inv_2 _0686_ (.A(_0111_),
    .Y(_0471_));
 sky130_fd_sc_hd__buf_8 _0687_ (.A(_0108_),
    .X(_0112_));
 sky130_fd_sc_hd__inv_2 _0688_ (.A(_0112_),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(_0112_),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(_0112_),
    .Y(_0474_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(_0112_),
    .Y(_0475_));
 sky130_fd_sc_hd__inv_2 _0692_ (.A(_0112_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _0693_ (.A(_0112_),
    .Y(_0477_));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(_0112_),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(_0112_),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(_0112_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _0697_ (.A(_0112_),
    .Y(_0487_));
 sky130_fd_sc_hd__buf_8 _0698_ (.A(_0108_),
    .X(_0113_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(_0113_),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(_0113_),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(_0113_),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_2 _0702_ (.A(_0113_),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(_0113_),
    .Y(_0481_));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(_0113_),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(_0113_),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(_0113_),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_2 _0707_ (.A(_0113_),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(_0113_),
    .Y(_0493_));
 sky130_fd_sc_hd__buf_12 _0709_ (.A(_0108_),
    .X(_0114_));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(_0114_),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(_0114_),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _0712_ (.A(_0114_),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(_0114_),
    .Y(_0497_));
 sky130_fd_sc_hd__inv_2 _0714_ (.A(_0114_),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(_0114_),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(_0114_),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(_0114_),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(_0114_),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _0719_ (.A(_0114_),
    .Y(_0503_));
 sky130_fd_sc_hd__buf_8 _0720_ (.A(_0108_),
    .X(_0115_));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(_0115_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(_0115_),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _0723_ (.A(_0115_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _0724_ (.A(_0115_),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_2 _0725_ (.A(_0115_),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(_0115_),
    .Y(_0509_));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(_0115_),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(_0115_),
    .Y(_0508_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(_0115_),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(_0115_),
    .Y(_0507_));
 sky130_fd_sc_hd__buf_8 _0731_ (.A(_0108_),
    .X(_0116_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(_0116_),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(_0116_),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(_0116_),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(_0116_),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(_0116_),
    .Y(_0519_));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(_0116_),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _0738_ (.A(_0116_),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(_0116_),
    .Y(_0523_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(_0116_),
    .Y(_0529_));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(_0116_),
    .Y(_0528_));
 sky130_fd_sc_hd__buf_8 _0742_ (.A(_0108_),
    .X(_0117_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(_0117_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(_0117_),
    .Y(_0527_));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(_0117_),
    .Y(_0531_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(_0117_),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_2 _0747_ (.A(_0117_),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(_0117_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(_0117_),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(_0117_),
    .Y(_0534_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(_0117_),
    .Y(_0535_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(_0117_),
    .Y(_0536_));
 sky130_fd_sc_hd__buf_8 _0753_ (.A(_0108_),
    .X(_0118_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(_0118_),
    .Y(_0537_));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(_0118_),
    .Y(_0538_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(_0118_),
    .Y(_0539_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(_0118_),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(_0118_),
    .Y(_0546_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(_0118_),
    .Y(_0545_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(_0118_),
    .Y(_0547_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(_0118_),
    .Y(_0544_));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(_0118_),
    .Y(_0548_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(_0118_),
    .Y(_0543_));
 sky130_fd_sc_hd__buf_8 _0764_ (.A(_0108_),
    .X(_0119_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(_0119_),
    .Y(_0549_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(_0119_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(_0119_),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(_0119_),
    .Y(_0551_));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(_0119_),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(_0119_),
    .Y(_0553_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(_0119_),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(_0119_),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(_0119_),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(_0119_),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(_0109_),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(_0109_),
    .Y(_0479_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(_0109_),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(_0109_),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(_0109_),
    .Y(_0541_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(_0109_),
    .Y(_0558_));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(_0109_),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(_0109_),
    .Y(_0483_));
 sky130_fd_sc_hd__inv_2 _0783_ (.A(\rgb_mixer.enc2[7] ),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(\rgb_mixer.enc2[6] ),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(\rgb_mixer.enc2[5] ),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(\rgb_mixer.enc2[4] ),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(\rgb_mixer.enc2[3] ),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(\rgb_mixer.enc2[2] ),
    .Y(_0125_));
 sky130_fd_sc_hd__o22a_1 _0789_ (.A1(_0124_),
    .A2(\rgb_mixer.pwm2.count[3] ),
    .B1(\rgb_mixer.pwm2.count[2] ),
    .B2(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(\rgb_mixer.enc2[0] ),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(\rgb_mixer.pwm2.count[7] ),
    .Y(_0128_));
 sky130_fd_sc_hd__a211o_1 _0792_ (.A1(_0127_),
    .A2(\rgb_mixer.pwm2.count[0] ),
    .B1(_0128_),
    .C1(\rgb_mixer.enc2[7] ),
    .X(_0129_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(\rgb_mixer.enc2[1] ),
    .Y(_0130_));
 sky130_fd_sc_hd__o22a_1 _0794_ (.A1(_0127_),
    .A2(\rgb_mixer.pwm2.count[0] ),
    .B1(\rgb_mixer.pwm2.count[1] ),
    .B2(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _0795_ (.A1(_0125_),
    .A2(\rgb_mixer.pwm2.count[2] ),
    .B1(\rgb_mixer.pwm2.count[1] ),
    .B2(_0130_),
    .X(_0132_));
 sky130_fd_sc_hd__a21o_1 _0796_ (.A1(_0129_),
    .A2(_0131_),
    .B1(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(_0123_),
    .A2(\rgb_mixer.pwm2.count[4] ),
    .B1(\rgb_mixer.pwm2.count[3] ),
    .B2(_0124_),
    .X(_0134_));
 sky130_fd_sc_hd__a21o_1 _0798_ (.A1(_0126_),
    .A2(_0133_),
    .B1(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__o221a_1 _0799_ (.A1(_0122_),
    .A2(\rgb_mixer.pwm2.count[5] ),
    .B1(\rgb_mixer.pwm2.count[4] ),
    .B2(_0123_),
    .C1(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__a221o_1 _0800_ (.A1(_0121_),
    .A2(\rgb_mixer.pwm2.count[6] ),
    .B1(\rgb_mixer.pwm2.count[5] ),
    .B2(_0122_),
    .C1(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__o221a_1 _0801_ (.A1(_0120_),
    .A2(\rgb_mixer.pwm2.count[7] ),
    .B1(\rgb_mixer.pwm2.count[6] ),
    .B2(_0121_),
    .C1(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_4 _0802_ (.A(net8),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_4 _0803_ (.A(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__a211oi_1 _0804_ (.A1(_0120_),
    .A2(\rgb_mixer.pwm2.count[7] ),
    .B1(_0138_),
    .C1(_0140_),
    .Y(\rgb_mixer.pwm2.out ));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(\rgb_mixer.enc1[7] ),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _0806_ (.A(\rgb_mixer.enc1[6] ),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _0807_ (.A(\rgb_mixer.enc1[5] ),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(\rgb_mixer.enc1[4] ),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(\rgb_mixer.enc1[3] ),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _0810_ (.A(\rgb_mixer.enc1[2] ),
    .Y(_0146_));
 sky130_fd_sc_hd__o22a_1 _0811_ (.A1(_0145_),
    .A2(\rgb_mixer.pwm1.count[3] ),
    .B1(\rgb_mixer.pwm1.count[2] ),
    .B2(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__inv_2 _0812_ (.A(\rgb_mixer.enc1[1] ),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(\rgb_mixer.enc1[0] ),
    .Y(_0149_));
 sky130_fd_sc_hd__and2_1 _0814_ (.A(_0149_),
    .B(\rgb_mixer.pwm1.count[0] ),
    .X(_0150_));
 sky130_fd_sc_hd__o2bb2a_1 _0815_ (.A1_N(_0141_),
    .A2_N(\rgb_mixer.pwm1.count[7] ),
    .B1(\rgb_mixer.pwm1.count[0] ),
    .B2(_0149_),
    .X(_0151_));
 sky130_fd_sc_hd__o22a_1 _0816_ (.A1(_0148_),
    .A2(\rgb_mixer.pwm1.count[1] ),
    .B1(_0150_),
    .B2(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__a221o_1 _0817_ (.A1(_0146_),
    .A2(\rgb_mixer.pwm1.count[2] ),
    .B1(\rgb_mixer.pwm1.count[1] ),
    .B2(_0148_),
    .C1(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _0818_ (.A(_0144_),
    .B(\rgb_mixer.pwm1.count[4] ),
    .X(_0154_));
 sky130_fd_sc_hd__a221o_1 _0819_ (.A1(_0145_),
    .A2(\rgb_mixer.pwm1.count[3] ),
    .B1(_0147_),
    .B2(_0153_),
    .C1(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__o221a_1 _0820_ (.A1(_0143_),
    .A2(\rgb_mixer.pwm1.count[5] ),
    .B1(\rgb_mixer.pwm1.count[4] ),
    .B2(_0144_),
    .C1(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__a221o_1 _0821_ (.A1(_0142_),
    .A2(\rgb_mixer.pwm1.count[6] ),
    .B1(\rgb_mixer.pwm1.count[5] ),
    .B2(_0143_),
    .C1(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__o22a_1 _0822_ (.A1(_0141_),
    .A2(\rgb_mixer.pwm1.count[7] ),
    .B1(\rgb_mixer.pwm1.count[6] ),
    .B2(_0142_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_4 _0823_ (.A(_0139_),
    .X(_0159_));
 sky130_fd_sc_hd__a221oi_1 _0824_ (.A1(_0141_),
    .A2(\rgb_mixer.pwm1.count[7] ),
    .B1(_0157_),
    .B2(_0158_),
    .C1(_0159_),
    .Y(\rgb_mixer.pwm1.out ));
 sky130_fd_sc_hd__inv_2 _0825_ (.A(_0139_),
    .Y(_0160_));
 sky130_fd_sc_hd__buf_2 _0826_ (.A(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_2 _0827_ (.A(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__or2b_1 _0828_ (.A(\rgb_mixer.enc0[7] ),
    .B_N(\rgb_mixer.pwm0.count[7] ),
    .X(_0163_));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(\rgb_mixer.pwm0.count[7] ),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(\rgb_mixer.pwm0.count[6] ),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _0831_ (.A(\rgb_mixer.pwm0.count[5] ),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(\rgb_mixer.pwm0.count[4] ),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(\rgb_mixer.pwm0.count[3] ),
    .Y(_0168_));
 sky130_fd_sc_hd__o22a_1 _0834_ (.A1(\rgb_mixer.enc0[4] ),
    .A2(_0167_),
    .B1(_0168_),
    .B2(\rgb_mixer.enc0[3] ),
    .X(_0169_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(\rgb_mixer.pwm0.count[2] ),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(\rgb_mixer.pwm0.count[1] ),
    .Y(_0171_));
 sky130_fd_sc_hd__o22a_1 _0837_ (.A1(\rgb_mixer.enc0[2] ),
    .A2(_0170_),
    .B1(_0171_),
    .B2(\rgb_mixer.enc0[1] ),
    .X(_0172_));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(\rgb_mixer.enc0[0] ),
    .Y(_0173_));
 sky130_fd_sc_hd__nand2_1 _0839_ (.A(_0173_),
    .B(\rgb_mixer.pwm0.count[0] ),
    .Y(_0174_));
 sky130_fd_sc_hd__o21ai_1 _0840_ (.A1(_0173_),
    .A2(\rgb_mixer.pwm0.count[0] ),
    .B1(_0163_),
    .Y(_0175_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(\rgb_mixer.enc0[1] ),
    .A2(_0171_),
    .B1(_0174_),
    .B2(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_1 _0842_ (.A1(\rgb_mixer.enc0[3] ),
    .A2(_0168_),
    .B1(_0170_),
    .B2(\rgb_mixer.enc0[2] ),
    .X(_0177_));
 sky130_fd_sc_hd__a21o_1 _0843_ (.A1(_0172_),
    .A2(_0176_),
    .B1(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_1 _0844_ (.A1(\rgb_mixer.enc0[5] ),
    .A2(_0166_),
    .B1(_0167_),
    .B2(\rgb_mixer.enc0[4] ),
    .X(_0179_));
 sky130_fd_sc_hd__a21o_1 _0845_ (.A1(_0169_),
    .A2(_0178_),
    .B1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__o221a_1 _0846_ (.A1(\rgb_mixer.enc0[6] ),
    .A2(_0165_),
    .B1(_0166_),
    .B2(\rgb_mixer.enc0[5] ),
    .C1(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__a221o_1 _0847_ (.A1(\rgb_mixer.enc0[7] ),
    .A2(_0164_),
    .B1(_0165_),
    .B2(\rgb_mixer.enc0[6] ),
    .C1(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__and3_1 _0848_ (.A(_0162_),
    .B(_0163_),
    .C(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _0849_ (.A(_0183_),
    .X(\rgb_mixer.pwm0.out ));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(\rgb_mixer.pwm2.count[0] ),
    .B(_0140_),
    .Y(_0000_));
 sky130_fd_sc_hd__a21oi_1 _0851_ (.A1(\rgb_mixer.pwm2.count[0] ),
    .A2(\rgb_mixer.pwm2.count[1] ),
    .B1(_0159_),
    .Y(_0184_));
 sky130_fd_sc_hd__o21a_1 _0852_ (.A1(\rgb_mixer.pwm2.count[0] ),
    .A2(\rgb_mixer.pwm2.count[1] ),
    .B1(_0184_),
    .X(_0001_));
 sky130_fd_sc_hd__a21oi_1 _0853_ (.A1(\rgb_mixer.pwm2.count[0] ),
    .A2(\rgb_mixer.pwm2.count[1] ),
    .B1(\rgb_mixer.pwm2.count[2] ),
    .Y(_0185_));
 sky130_fd_sc_hd__and3_1 _0854_ (.A(\rgb_mixer.pwm2.count[0] ),
    .B(\rgb_mixer.pwm2.count[2] ),
    .C(\rgb_mixer.pwm2.count[1] ),
    .X(_0186_));
 sky130_fd_sc_hd__nor3_1 _0855_ (.A(_0140_),
    .B(_0185_),
    .C(_0186_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2_1 _0856_ (.A(\rgb_mixer.pwm2.count[3] ),
    .B(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_4 _0857_ (.A(_0161_),
    .X(_0188_));
 sky130_fd_sc_hd__o21ai_1 _0858_ (.A1(\rgb_mixer.pwm2.count[3] ),
    .A2(_0186_),
    .B1(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _0859_ (.A(_0187_),
    .B(_0189_),
    .Y(_0003_));
 sky130_fd_sc_hd__a21oi_1 _0860_ (.A1(\rgb_mixer.pwm2.count[4] ),
    .A2(_0187_),
    .B1(_0159_),
    .Y(_0190_));
 sky130_fd_sc_hd__o21a_1 _0861_ (.A1(\rgb_mixer.pwm2.count[4] ),
    .A2(_0187_),
    .B1(_0190_),
    .X(_0004_));
 sky130_fd_sc_hd__a21oi_1 _0862_ (.A1(\rgb_mixer.pwm2.count[4] ),
    .A2(_0187_),
    .B1(\rgb_mixer.pwm2.count[5] ),
    .Y(_0191_));
 sky130_fd_sc_hd__and3_1 _0863_ (.A(\rgb_mixer.pwm2.count[5] ),
    .B(\rgb_mixer.pwm2.count[4] ),
    .C(_0187_),
    .X(_0192_));
 sky130_fd_sc_hd__nor3_1 _0864_ (.A(_0140_),
    .B(_0191_),
    .C(_0192_),
    .Y(_0005_));
 sky130_fd_sc_hd__and2_1 _0865_ (.A(\rgb_mixer.pwm2.count[6] ),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__o21ai_1 _0866_ (.A1(\rgb_mixer.pwm2.count[6] ),
    .A2(_0192_),
    .B1(_0188_),
    .Y(_0194_));
 sky130_fd_sc_hd__nor2_1 _0867_ (.A(_0193_),
    .B(_0194_),
    .Y(_0006_));
 sky130_fd_sc_hd__a21oi_1 _0868_ (.A1(\rgb_mixer.pwm2.count[7] ),
    .A2(_0193_),
    .B1(_0159_),
    .Y(_0195_));
 sky130_fd_sc_hd__o21a_1 _0869_ (.A1(\rgb_mixer.pwm2.count[7] ),
    .A2(_0193_),
    .B1(_0195_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_1 _0870_ (.A(_0140_),
    .B(\rgb_mixer.pwm1.count[0] ),
    .Y(_0008_));
 sky130_fd_sc_hd__a21oi_1 _0871_ (.A1(\rgb_mixer.pwm1.count[1] ),
    .A2(\rgb_mixer.pwm1.count[0] ),
    .B1(_0159_),
    .Y(_0196_));
 sky130_fd_sc_hd__o21a_1 _0872_ (.A1(\rgb_mixer.pwm1.count[1] ),
    .A2(\rgb_mixer.pwm1.count[0] ),
    .B1(_0196_),
    .X(_0009_));
 sky130_fd_sc_hd__a21oi_1 _0873_ (.A1(\rgb_mixer.pwm1.count[1] ),
    .A2(\rgb_mixer.pwm1.count[0] ),
    .B1(\rgb_mixer.pwm1.count[2] ),
    .Y(_0197_));
 sky130_fd_sc_hd__and3_1 _0874_ (.A(\rgb_mixer.pwm1.count[2] ),
    .B(\rgb_mixer.pwm1.count[1] ),
    .C(\rgb_mixer.pwm1.count[0] ),
    .X(_0198_));
 sky130_fd_sc_hd__nor3_1 _0875_ (.A(_0140_),
    .B(_0197_),
    .C(_0198_),
    .Y(_0010_));
 sky130_fd_sc_hd__and2_1 _0876_ (.A(\rgb_mixer.pwm1.count[3] ),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__o21ai_1 _0877_ (.A1(\rgb_mixer.pwm1.count[3] ),
    .A2(_0198_),
    .B1(_0188_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _0878_ (.A(_0199_),
    .B(_0200_),
    .Y(_0011_));
 sky130_fd_sc_hd__and3_1 _0879_ (.A(\rgb_mixer.pwm1.count[4] ),
    .B(\rgb_mixer.pwm1.count[3] ),
    .C(_0198_),
    .X(_0201_));
 sky130_fd_sc_hd__o21ai_1 _0880_ (.A1(\rgb_mixer.pwm1.count[4] ),
    .A2(_0199_),
    .B1(_0188_),
    .Y(_0202_));
 sky130_fd_sc_hd__nor2_1 _0881_ (.A(_0201_),
    .B(_0202_),
    .Y(_0012_));
 sky130_fd_sc_hd__and2_1 _0882_ (.A(\rgb_mixer.pwm1.count[5] ),
    .B(_0201_),
    .X(_0203_));
 sky130_fd_sc_hd__nor2_1 _0883_ (.A(_0139_),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__o21a_1 _0884_ (.A1(\rgb_mixer.pwm1.count[5] ),
    .A2(_0201_),
    .B1(_0204_),
    .X(_0013_));
 sky130_fd_sc_hd__and3_1 _0885_ (.A(\rgb_mixer.pwm1.count[6] ),
    .B(\rgb_mixer.pwm1.count[5] ),
    .C(_0201_),
    .X(_0205_));
 sky130_fd_sc_hd__o21ai_1 _0886_ (.A1(\rgb_mixer.pwm1.count[6] ),
    .A2(_0203_),
    .B1(_0188_),
    .Y(_0206_));
 sky130_fd_sc_hd__nor2_1 _0887_ (.A(_0205_),
    .B(_0206_),
    .Y(_0014_));
 sky130_fd_sc_hd__a21oi_1 _0888_ (.A1(\rgb_mixer.pwm1.count[7] ),
    .A2(_0205_),
    .B1(_0159_),
    .Y(_0207_));
 sky130_fd_sc_hd__o21a_1 _0889_ (.A1(\rgb_mixer.pwm1.count[7] ),
    .A2(_0205_),
    .B1(_0207_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_1 _0890_ (.A(_0140_),
    .B(\rgb_mixer.pwm0.count[0] ),
    .Y(_0016_));
 sky130_fd_sc_hd__a21oi_1 _0891_ (.A1(\rgb_mixer.pwm0.count[1] ),
    .A2(\rgb_mixer.pwm0.count[0] ),
    .B1(_0159_),
    .Y(_0208_));
 sky130_fd_sc_hd__o21a_1 _0892_ (.A1(\rgb_mixer.pwm0.count[1] ),
    .A2(\rgb_mixer.pwm0.count[0] ),
    .B1(_0208_),
    .X(_0017_));
 sky130_fd_sc_hd__a21oi_1 _0893_ (.A1(\rgb_mixer.pwm0.count[1] ),
    .A2(\rgb_mixer.pwm0.count[0] ),
    .B1(\rgb_mixer.pwm0.count[2] ),
    .Y(_0209_));
 sky130_fd_sc_hd__and3_1 _0894_ (.A(\rgb_mixer.pwm0.count[2] ),
    .B(\rgb_mixer.pwm0.count[1] ),
    .C(\rgb_mixer.pwm0.count[0] ),
    .X(_0210_));
 sky130_fd_sc_hd__nor3_1 _0895_ (.A(_0140_),
    .B(_0209_),
    .C(_0210_),
    .Y(_0018_));
 sky130_fd_sc_hd__and2_1 _0896_ (.A(\rgb_mixer.pwm0.count[3] ),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__o21ai_1 _0897_ (.A1(\rgb_mixer.pwm0.count[3] ),
    .A2(_0210_),
    .B1(_0188_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _0898_ (.A(_0211_),
    .B(_0212_),
    .Y(_0019_));
 sky130_fd_sc_hd__a21oi_1 _0899_ (.A1(\rgb_mixer.pwm0.count[4] ),
    .A2(_0211_),
    .B1(_0139_),
    .Y(_0213_));
 sky130_fd_sc_hd__o21a_1 _0900_ (.A1(\rgb_mixer.pwm0.count[4] ),
    .A2(_0211_),
    .B1(_0213_),
    .X(_0020_));
 sky130_fd_sc_hd__a21oi_1 _0901_ (.A1(\rgb_mixer.pwm0.count[4] ),
    .A2(_0211_),
    .B1(\rgb_mixer.pwm0.count[5] ),
    .Y(_0214_));
 sky130_fd_sc_hd__and3_1 _0902_ (.A(\rgb_mixer.pwm0.count[5] ),
    .B(\rgb_mixer.pwm0.count[4] ),
    .C(_0211_),
    .X(_0215_));
 sky130_fd_sc_hd__nor3_1 _0903_ (.A(_0140_),
    .B(_0214_),
    .C(_0215_),
    .Y(_0021_));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(\rgb_mixer.pwm0.count[6] ),
    .B(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__o21ai_1 _0905_ (.A1(\rgb_mixer.pwm0.count[6] ),
    .A2(_0215_),
    .B1(_0188_),
    .Y(_0217_));
 sky130_fd_sc_hd__nor2_1 _0906_ (.A(_0216_),
    .B(_0217_),
    .Y(_0022_));
 sky130_fd_sc_hd__a21oi_1 _0907_ (.A1(\rgb_mixer.pwm0.count[7] ),
    .A2(_0216_),
    .B1(_0139_),
    .Y(_0218_));
 sky130_fd_sc_hd__o21a_1 _0908_ (.A1(\rgb_mixer.pwm0.count[7] ),
    .A2(_0216_),
    .B1(_0218_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _0909_ (.A(\rgb_mixer.debounce2_b.debounced ),
    .B(_0161_),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_1 _0910_ (.A(_0219_),
    .X(_0024_));
 sky130_fd_sc_hd__and2b_1 _0911_ (.A_N(\rgb_mixer.debounce2_a.debounced ),
    .B(\rgb_mixer.debounce2_b.debounced ),
    .X(_0220_));
 sky130_fd_sc_hd__and2b_1 _0912_ (.A_N(\rgb_mixer.debounce2_b.debounced ),
    .B(\rgb_mixer.debounce2_a.debounced ),
    .X(_0221_));
 sky130_fd_sc_hd__and2_1 _0913_ (.A(\rgb_mixer.encoder2.old_b ),
    .B(\rgb_mixer.encoder2.old_a ),
    .X(_0222_));
 sky130_fd_sc_hd__nor2_1 _0914_ (.A(\rgb_mixer.encoder2.old_b ),
    .B(\rgb_mixer.encoder2.old_a ),
    .Y(_0223_));
 sky130_fd_sc_hd__o22a_2 _0915_ (.A1(_0220_),
    .A2(_0221_),
    .B1(_0222_),
    .B2(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_4 _0916_ (.A(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__a21oi_1 _0917_ (.A1(\rgb_mixer.enc2[0] ),
    .A2(_0224_),
    .B1(_0139_),
    .Y(_0226_));
 sky130_fd_sc_hd__o21a_1 _0918_ (.A1(\rgb_mixer.enc2[0] ),
    .A2(_0225_),
    .B1(_0226_),
    .X(_0025_));
 sky130_fd_sc_hd__and4b_1 _0919_ (.A_N(\rgb_mixer.debounce2_b.debounced ),
    .B(\rgb_mixer.encoder2.old_b ),
    .C(\rgb_mixer.encoder2.old_a ),
    .D(\rgb_mixer.debounce2_a.debounced ),
    .X(_0227_));
 sky130_fd_sc_hd__a21o_1 _0920_ (.A1(_0220_),
    .A2(_0223_),
    .B1(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_4 _0921_ (.A(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__nor2_1 _0922_ (.A(\rgb_mixer.enc2[1] ),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__o221a_1 _0923_ (.A1(_0220_),
    .A2(_0222_),
    .B1(_0223_),
    .B2(_0221_),
    .C1(\rgb_mixer.enc2[1] ),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _0924_ (.A(_0230_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__xnor2_1 _0925_ (.A(\rgb_mixer.enc2[0] ),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _0926_ (.A(_0225_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__buf_4 _0927_ (.A(_0162_),
    .X(_0235_));
 sky130_fd_sc_hd__o211a_1 _0928_ (.A1(\rgb_mixer.enc2[1] ),
    .A2(_0225_),
    .B1(_0234_),
    .C1(_0235_),
    .X(_0026_));
 sky130_fd_sc_hd__a211o_1 _0929_ (.A1(_0220_),
    .A2(_0223_),
    .B1(_0227_),
    .C1(\rgb_mixer.enc2[1] ),
    .X(_0236_));
 sky130_fd_sc_hd__a21o_1 _0930_ (.A1(\rgb_mixer.enc2[0] ),
    .A2(_0236_),
    .B1(_0231_),
    .X(_0237_));
 sky130_fd_sc_hd__xnor2_1 _0931_ (.A(_0125_),
    .B(_0228_),
    .Y(_0238_));
 sky130_fd_sc_hd__or2_1 _0932_ (.A(_0237_),
    .B(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _0933_ (.A(_0237_),
    .B(_0238_),
    .Y(_0240_));
 sky130_fd_sc_hd__a21bo_1 _0934_ (.A1(_0239_),
    .A2(_0240_),
    .B1_N(_0224_),
    .X(_0241_));
 sky130_fd_sc_hd__o211a_1 _0935_ (.A1(\rgb_mixer.enc2[2] ),
    .A2(_0225_),
    .B1(_0241_),
    .C1(_0235_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _0936_ (.A(\rgb_mixer.enc2[2] ),
    .B(_0229_),
    .Y(_0242_));
 sky130_fd_sc_hd__xnor2_1 _0937_ (.A(_0124_),
    .B(_0228_),
    .Y(_0243_));
 sky130_fd_sc_hd__and3_1 _0938_ (.A(_0242_),
    .B(_0240_),
    .C(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__a21o_1 _0939_ (.A1(_0242_),
    .A2(_0240_),
    .B1(_0243_),
    .X(_0245_));
 sky130_fd_sc_hd__nand2_1 _0940_ (.A(_0224_),
    .B(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__buf_4 _0941_ (.A(_0161_),
    .X(_0247_));
 sky130_fd_sc_hd__o221a_1 _0942_ (.A1(\rgb_mixer.enc2[3] ),
    .A2(_0225_),
    .B1(_0244_),
    .B2(_0246_),
    .C1(_0247_),
    .X(_0028_));
 sky130_fd_sc_hd__o21a_1 _0943_ (.A1(\rgb_mixer.enc2[3] ),
    .A2(\rgb_mixer.enc2[2] ),
    .B1(_0229_),
    .X(_0248_));
 sky130_fd_sc_hd__a31o_1 _0944_ (.A1(_0237_),
    .A2(_0238_),
    .A3(_0243_),
    .B1(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__xnor2_1 _0945_ (.A(_0123_),
    .B(_0229_),
    .Y(_0250_));
 sky130_fd_sc_hd__or2_1 _0946_ (.A(_0249_),
    .B(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _0947_ (.A(_0249_),
    .B(_0250_),
    .Y(_0252_));
 sky130_fd_sc_hd__a21bo_1 _0948_ (.A1(_0251_),
    .A2(_0252_),
    .B1_N(_0224_),
    .X(_0253_));
 sky130_fd_sc_hd__o211a_1 _0949_ (.A1(\rgb_mixer.enc2[4] ),
    .A2(_0225_),
    .B1(_0253_),
    .C1(_0235_),
    .X(_0029_));
 sky130_fd_sc_hd__xnor2_1 _0950_ (.A(_0122_),
    .B(_0229_),
    .Y(_0254_));
 sky130_fd_sc_hd__a21bo_1 _0951_ (.A1(\rgb_mixer.enc2[4] ),
    .A2(_0229_),
    .B1_N(_0252_),
    .X(_0255_));
 sky130_fd_sc_hd__xnor2_1 _0952_ (.A(_0254_),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor2_1 _0953_ (.A(\rgb_mixer.enc2[5] ),
    .B(_0224_),
    .Y(_0257_));
 sky130_fd_sc_hd__a211oi_1 _0954_ (.A1(_0225_),
    .A2(_0256_),
    .B1(_0257_),
    .C1(_0140_),
    .Y(_0030_));
 sky130_fd_sc_hd__nor2_1 _0955_ (.A(\rgb_mixer.enc2[6] ),
    .B(_0229_),
    .Y(_0258_));
 sky130_fd_sc_hd__and2_1 _0956_ (.A(\rgb_mixer.enc2[6] ),
    .B(_0229_),
    .X(_0259_));
 sky130_fd_sc_hd__nor2_1 _0957_ (.A(_0258_),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__o21a_1 _0958_ (.A1(\rgb_mixer.enc2[5] ),
    .A2(\rgb_mixer.enc2[4] ),
    .B1(_0229_),
    .X(_0261_));
 sky130_fd_sc_hd__a31o_1 _0959_ (.A1(_0249_),
    .A2(_0250_),
    .A3(_0254_),
    .B1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__xnor2_1 _0960_ (.A(_0260_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _0961_ (.A(_0225_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__o211a_1 _0962_ (.A1(\rgb_mixer.enc2[6] ),
    .A2(_0225_),
    .B1(_0264_),
    .C1(_0235_),
    .X(_0031_));
 sky130_fd_sc_hd__a21o_1 _0963_ (.A1(_0260_),
    .A2(_0262_),
    .B1(_0259_),
    .X(_0265_));
 sky130_fd_sc_hd__xnor2_1 _0964_ (.A(_0120_),
    .B(_0229_),
    .Y(_0266_));
 sky130_fd_sc_hd__xnor2_1 _0965_ (.A(_0265_),
    .B(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__nor2_1 _0966_ (.A(\rgb_mixer.enc2[7] ),
    .B(_0224_),
    .Y(_0268_));
 sky130_fd_sc_hd__a211oi_1 _0967_ (.A1(_0225_),
    .A2(_0267_),
    .B1(_0268_),
    .C1(_0159_),
    .Y(_0032_));
 sky130_fd_sc_hd__clkbuf_4 _0968_ (.A(_0161_),
    .X(_0269_));
 sky130_fd_sc_hd__and2_1 _0969_ (.A(\rgb_mixer.debounce1_b.debounced ),
    .B(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _0970_ (.A(_0270_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _0971_ (.A(\rgb_mixer.debounce2_a.debounced ),
    .B(_0269_),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _0972_ (.A(_0271_),
    .X(_0034_));
 sky130_fd_sc_hd__and2b_1 _0973_ (.A_N(\rgb_mixer.debounce1_a.debounced ),
    .B(\rgb_mixer.debounce1_b.debounced ),
    .X(_0272_));
 sky130_fd_sc_hd__and2b_1 _0974_ (.A_N(\rgb_mixer.debounce1_b.debounced ),
    .B(\rgb_mixer.debounce1_a.debounced ),
    .X(_0273_));
 sky130_fd_sc_hd__and2_1 _0975_ (.A(\rgb_mixer.encoder1.old_b ),
    .B(\rgb_mixer.encoder1.old_a ),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_1 _0976_ (.A(\rgb_mixer.encoder1.old_b ),
    .B(\rgb_mixer.encoder1.old_a ),
    .Y(_0275_));
 sky130_fd_sc_hd__o22a_2 _0977_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0274_),
    .B2(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__buf_2 _0978_ (.A(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__a21oi_1 _0979_ (.A1(\rgb_mixer.enc1[0] ),
    .A2(_0276_),
    .B1(_0139_),
    .Y(_0278_));
 sky130_fd_sc_hd__o21a_1 _0980_ (.A1(\rgb_mixer.enc1[0] ),
    .A2(_0277_),
    .B1(_0278_),
    .X(_0035_));
 sky130_fd_sc_hd__and4b_1 _0981_ (.A_N(\rgb_mixer.debounce1_b.debounced ),
    .B(\rgb_mixer.encoder1.old_b ),
    .C(\rgb_mixer.encoder1.old_a ),
    .D(\rgb_mixer.debounce1_a.debounced ),
    .X(_0279_));
 sky130_fd_sc_hd__a21o_1 _0982_ (.A1(_0272_),
    .A2(_0275_),
    .B1(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_4 _0983_ (.A(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__nor2_1 _0984_ (.A(\rgb_mixer.enc1[1] ),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__o221a_1 _0985_ (.A1(_0272_),
    .A2(_0274_),
    .B1(_0275_),
    .B2(_0273_),
    .C1(\rgb_mixer.enc1[1] ),
    .X(_0283_));
 sky130_fd_sc_hd__nor2_1 _0986_ (.A(_0282_),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__xnor2_1 _0987_ (.A(\rgb_mixer.enc1[0] ),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand2_1 _0988_ (.A(_0277_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__o211a_1 _0989_ (.A1(\rgb_mixer.enc1[1] ),
    .A2(_0277_),
    .B1(_0286_),
    .C1(_0235_),
    .X(_0036_));
 sky130_fd_sc_hd__a211o_1 _0990_ (.A1(_0272_),
    .A2(_0275_),
    .B1(_0279_),
    .C1(\rgb_mixer.enc1[1] ),
    .X(_0287_));
 sky130_fd_sc_hd__a21o_1 _0991_ (.A1(\rgb_mixer.enc1[0] ),
    .A2(_0287_),
    .B1(_0283_),
    .X(_0288_));
 sky130_fd_sc_hd__xnor2_1 _0992_ (.A(_0146_),
    .B(_0280_),
    .Y(_0289_));
 sky130_fd_sc_hd__or2_1 _0993_ (.A(_0288_),
    .B(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__nand2_1 _0994_ (.A(_0288_),
    .B(_0289_),
    .Y(_0291_));
 sky130_fd_sc_hd__a21bo_1 _0995_ (.A1(_0290_),
    .A2(_0291_),
    .B1_N(_0276_),
    .X(_0292_));
 sky130_fd_sc_hd__o211a_1 _0996_ (.A1(\rgb_mixer.enc1[2] ),
    .A2(_0277_),
    .B1(_0292_),
    .C1(_0235_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _0997_ (.A(\rgb_mixer.enc1[2] ),
    .B(_0281_),
    .Y(_0293_));
 sky130_fd_sc_hd__xnor2_1 _0998_ (.A(_0145_),
    .B(_0280_),
    .Y(_0294_));
 sky130_fd_sc_hd__and3_1 _0999_ (.A(_0293_),
    .B(_0291_),
    .C(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__a21o_1 _1000_ (.A1(_0293_),
    .A2(_0291_),
    .B1(_0294_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(_0276_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__o221a_1 _1002_ (.A1(\rgb_mixer.enc1[3] ),
    .A2(_0277_),
    .B1(_0295_),
    .B2(_0297_),
    .C1(_0247_),
    .X(_0038_));
 sky130_fd_sc_hd__o21a_1 _1003_ (.A1(\rgb_mixer.enc1[3] ),
    .A2(\rgb_mixer.enc1[2] ),
    .B1(_0281_),
    .X(_0298_));
 sky130_fd_sc_hd__a31o_1 _1004_ (.A1(_0288_),
    .A2(_0289_),
    .A3(_0294_),
    .B1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__xnor2_1 _1005_ (.A(_0144_),
    .B(_0281_),
    .Y(_0300_));
 sky130_fd_sc_hd__or2_1 _1006_ (.A(_0299_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(_0299_),
    .B(_0300_),
    .Y(_0302_));
 sky130_fd_sc_hd__a21bo_1 _1008_ (.A1(_0301_),
    .A2(_0302_),
    .B1_N(_0276_),
    .X(_0303_));
 sky130_fd_sc_hd__o211a_1 _1009_ (.A1(\rgb_mixer.enc1[4] ),
    .A2(_0277_),
    .B1(_0303_),
    .C1(_0235_),
    .X(_0039_));
 sky130_fd_sc_hd__xnor2_1 _1010_ (.A(_0143_),
    .B(_0281_),
    .Y(_0304_));
 sky130_fd_sc_hd__a21bo_1 _1011_ (.A1(\rgb_mixer.enc1[4] ),
    .A2(_0281_),
    .B1_N(_0302_),
    .X(_0305_));
 sky130_fd_sc_hd__xnor2_1 _1012_ (.A(_0304_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(\rgb_mixer.enc1[5] ),
    .B(_0276_),
    .Y(_0307_));
 sky130_fd_sc_hd__a211oi_1 _1014_ (.A1(_0277_),
    .A2(_0306_),
    .B1(_0307_),
    .C1(_0159_),
    .Y(_0040_));
 sky130_fd_sc_hd__nor2_1 _1015_ (.A(\rgb_mixer.enc1[6] ),
    .B(_0281_),
    .Y(_0308_));
 sky130_fd_sc_hd__and2_1 _1016_ (.A(\rgb_mixer.enc1[6] ),
    .B(_0281_),
    .X(_0309_));
 sky130_fd_sc_hd__nor2_1 _1017_ (.A(_0308_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__o21a_1 _1018_ (.A1(\rgb_mixer.enc1[5] ),
    .A2(\rgb_mixer.enc1[4] ),
    .B1(_0281_),
    .X(_0311_));
 sky130_fd_sc_hd__a31o_1 _1019_ (.A1(_0299_),
    .A2(_0300_),
    .A3(_0304_),
    .B1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__xnor2_1 _1020_ (.A(_0310_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _1021_ (.A(_0277_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__o211a_1 _1022_ (.A1(\rgb_mixer.enc1[6] ),
    .A2(_0277_),
    .B1(_0314_),
    .C1(_0235_),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _1023_ (.A1(_0310_),
    .A2(_0312_),
    .B1(_0309_),
    .X(_0315_));
 sky130_fd_sc_hd__xnor2_1 _1024_ (.A(_0141_),
    .B(_0281_),
    .Y(_0316_));
 sky130_fd_sc_hd__xnor2_1 _1025_ (.A(_0315_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nor2_1 _1026_ (.A(\rgb_mixer.enc1[7] ),
    .B(_0276_),
    .Y(_0318_));
 sky130_fd_sc_hd__a211oi_1 _1027_ (.A1(_0277_),
    .A2(_0317_),
    .B1(_0318_),
    .C1(_0159_),
    .Y(_0042_));
 sky130_fd_sc_hd__and2_1 _1028_ (.A(\rgb_mixer.debounce0_b.debounced ),
    .B(_0269_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _1029_ (.A(_0319_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _1030_ (.A(\rgb_mixer.debounce1_a.debounced ),
    .B(_0269_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0320_),
    .X(_0044_));
 sky130_fd_sc_hd__and2b_1 _1032_ (.A_N(\rgb_mixer.debounce0_a.debounced ),
    .B(\rgb_mixer.debounce0_b.debounced ),
    .X(_0321_));
 sky130_fd_sc_hd__and2b_1 _1033_ (.A_N(\rgb_mixer.debounce0_b.debounced ),
    .B(\rgb_mixer.debounce0_a.debounced ),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _1034_ (.A(\rgb_mixer.encoder0.old_b ),
    .B(\rgb_mixer.encoder0.old_a ),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_1 _1035_ (.A(\rgb_mixer.encoder0.old_b ),
    .B(\rgb_mixer.encoder0.old_a ),
    .Y(_0324_));
 sky130_fd_sc_hd__o22a_1 _1036_ (.A1(_0321_),
    .A2(_0322_),
    .B1(_0323_),
    .B2(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__clkinv_2 _1037_ (.A(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__buf_2 _1038_ (.A(_0325_),
    .X(_0327_));
 sky130_fd_sc_hd__a21o_1 _1039_ (.A1(\rgb_mixer.enc0[0] ),
    .A2(_0327_),
    .B1(_0139_),
    .X(_0328_));
 sky130_fd_sc_hd__a21oi_1 _1040_ (.A1(_0173_),
    .A2(_0326_),
    .B1(_0328_),
    .Y(_0045_));
 sky130_fd_sc_hd__and4b_1 _1041_ (.A_N(\rgb_mixer.debounce0_b.debounced ),
    .B(\rgb_mixer.encoder0.old_b ),
    .C(\rgb_mixer.encoder0.old_a ),
    .D(\rgb_mixer.debounce0_a.debounced ),
    .X(_0329_));
 sky130_fd_sc_hd__a21o_1 _1042_ (.A1(_0321_),
    .A2(_0324_),
    .B1(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_4 _1043_ (.A(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_1 _1044_ (.A(\rgb_mixer.enc0[1] ),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__o221a_1 _1045_ (.A1(_0321_),
    .A2(_0323_),
    .B1(_0324_),
    .B2(_0322_),
    .C1(\rgb_mixer.enc0[1] ),
    .X(_0333_));
 sky130_fd_sc_hd__nor2_1 _1046_ (.A(_0332_),
    .B(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__or2_1 _1047_ (.A(\rgb_mixer.enc0[0] ),
    .B(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(\rgb_mixer.enc0[0] ),
    .B(_0334_),
    .Y(_0336_));
 sky130_fd_sc_hd__a21o_1 _1049_ (.A1(_0335_),
    .A2(_0336_),
    .B1(_0326_),
    .X(_0337_));
 sky130_fd_sc_hd__o211a_1 _1050_ (.A1(\rgb_mixer.enc0[1] ),
    .A2(_0327_),
    .B1(_0337_),
    .C1(_0235_),
    .X(_0046_));
 sky130_fd_sc_hd__a211o_1 _1051_ (.A1(_0321_),
    .A2(_0324_),
    .B1(_0329_),
    .C1(\rgb_mixer.enc0[1] ),
    .X(_0338_));
 sky130_fd_sc_hd__a21o_1 _1052_ (.A1(\rgb_mixer.enc0[0] ),
    .A2(_0338_),
    .B1(_0333_),
    .X(_0339_));
 sky130_fd_sc_hd__xor2_1 _1053_ (.A(\rgb_mixer.enc0[2] ),
    .B(_0330_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _1054_ (.A(_0339_),
    .B(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(_0339_),
    .B(_0340_),
    .Y(_0342_));
 sky130_fd_sc_hd__a21o_1 _1056_ (.A1(_0341_),
    .A2(_0342_),
    .B1(_0326_),
    .X(_0343_));
 sky130_fd_sc_hd__o211a_1 _1057_ (.A1(\rgb_mixer.enc0[2] ),
    .A2(_0327_),
    .B1(_0343_),
    .C1(_0235_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _1058_ (.A(\rgb_mixer.enc0[2] ),
    .B(_0331_),
    .Y(_0344_));
 sky130_fd_sc_hd__xor2_1 _1059_ (.A(\rgb_mixer.enc0[3] ),
    .B(_0330_),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_1 _1060_ (.A1(_0344_),
    .A2(_0342_),
    .B1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a31o_1 _1061_ (.A1(_0344_),
    .A2(_0342_),
    .A3(_0345_),
    .B1(_0326_),
    .X(_0347_));
 sky130_fd_sc_hd__o221a_1 _1062_ (.A1(\rgb_mixer.enc0[3] ),
    .A2(_0327_),
    .B1(_0346_),
    .B2(_0347_),
    .C1(_0247_),
    .X(_0048_));
 sky130_fd_sc_hd__o21a_1 _1063_ (.A1(\rgb_mixer.enc0[3] ),
    .A2(\rgb_mixer.enc0[2] ),
    .B1(_0331_),
    .X(_0348_));
 sky130_fd_sc_hd__a31o_1 _1064_ (.A1(_0339_),
    .A2(_0340_),
    .A3(_0345_),
    .B1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__xor2_1 _1065_ (.A(\rgb_mixer.enc0[4] ),
    .B(_0331_),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _1066_ (.A(_0349_),
    .B(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _1067_ (.A(_0349_),
    .B(_0350_),
    .Y(_0352_));
 sky130_fd_sc_hd__a21o_1 _1068_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0326_),
    .X(_0353_));
 sky130_fd_sc_hd__o211a_1 _1069_ (.A1(\rgb_mixer.enc0[4] ),
    .A2(_0327_),
    .B1(_0353_),
    .C1(_0247_),
    .X(_0049_));
 sky130_fd_sc_hd__xor2_1 _1070_ (.A(\rgb_mixer.enc0[5] ),
    .B(_0331_),
    .X(_0354_));
 sky130_fd_sc_hd__a21bo_1 _1071_ (.A1(\rgb_mixer.enc0[4] ),
    .A2(_0331_),
    .B1_N(_0352_),
    .X(_0355_));
 sky130_fd_sc_hd__xnor2_1 _1072_ (.A(_0354_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__o21ai_1 _1073_ (.A1(\rgb_mixer.enc0[5] ),
    .A2(_0327_),
    .B1(_0188_),
    .Y(_0357_));
 sky130_fd_sc_hd__a21oi_1 _1074_ (.A1(_0327_),
    .A2(_0356_),
    .B1(_0357_),
    .Y(_0050_));
 sky130_fd_sc_hd__nor2_1 _1075_ (.A(\rgb_mixer.enc0[6] ),
    .B(_0331_),
    .Y(_0358_));
 sky130_fd_sc_hd__and2_1 _1076_ (.A(\rgb_mixer.enc0[6] ),
    .B(_0331_),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_1 _1077_ (.A(_0358_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__o21a_1 _1078_ (.A1(\rgb_mixer.enc0[5] ),
    .A2(\rgb_mixer.enc0[4] ),
    .B1(_0331_),
    .X(_0361_));
 sky130_fd_sc_hd__a31o_1 _1079_ (.A1(_0349_),
    .A2(_0350_),
    .A3(_0354_),
    .B1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__xor2_1 _1080_ (.A(_0360_),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _1081_ (.A(\rgb_mixer.enc0[6] ),
    .B(_0327_),
    .X(_0364_));
 sky130_fd_sc_hd__o211a_1 _1082_ (.A1(_0326_),
    .A2(_0363_),
    .B1(_0364_),
    .C1(_0247_),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _1083_ (.A1(_0360_),
    .A2(_0362_),
    .B1(_0359_),
    .X(_0365_));
 sky130_fd_sc_hd__xor2_1 _1084_ (.A(\rgb_mixer.enc0[7] ),
    .B(_0331_),
    .X(_0366_));
 sky130_fd_sc_hd__xnor2_1 _1085_ (.A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__o21ai_1 _1086_ (.A1(\rgb_mixer.enc0[7] ),
    .A2(_0327_),
    .B1(_0188_),
    .Y(_0368_));
 sky130_fd_sc_hd__a21oi_1 _1087_ (.A1(_0327_),
    .A2(_0367_),
    .B1(_0368_),
    .Y(_0052_));
 sky130_fd_sc_hd__and2_1 _1088_ (.A(_0269_),
    .B(net5),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _1089_ (.A(_0369_),
    .X(_0053_));
 sky130_fd_sc_hd__clkbuf_2 _1090_ (.A(_0161_),
    .X(_0370_));
 sky130_fd_sc_hd__and2_1 _1091_ (.A(\rgb_mixer.debounce2_b.button_hist[0] ),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _1092_ (.A(_0371_),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _1093_ (.A(\rgb_mixer.debounce2_b.button_hist[1] ),
    .B(_0370_),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _1094_ (.A(_0372_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _1095_ (.A(\rgb_mixer.debounce2_b.button_hist[2] ),
    .B(_0370_),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _1096_ (.A(_0373_),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _1097_ (.A(\rgb_mixer.debounce2_b.button_hist[3] ),
    .B(_0370_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _1098_ (.A(_0374_),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _1099_ (.A(\rgb_mixer.debounce2_b.button_hist[4] ),
    .B(_0370_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _1100_ (.A(_0375_),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _1101_ (.A(\rgb_mixer.debounce2_b.button_hist[5] ),
    .B(_0370_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _1102_ (.A(_0376_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _1103_ (.A(\rgb_mixer.debounce2_b.button_hist[6] ),
    .B(_0370_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _1104_ (.A(_0377_),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _1105_ (.A(\rgb_mixer.debounce0_a.debounced ),
    .B(_0161_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _1106_ (.A(_0378_),
    .X(_0061_));
 sky130_fd_sc_hd__and4_1 _1107_ (.A(\rgb_mixer.debounce2_b.button_hist[4] ),
    .B(\rgb_mixer.debounce2_b.button_hist[5] ),
    .C(\rgb_mixer.debounce2_b.button_hist[7] ),
    .D(\rgb_mixer.debounce2_b.button_hist[6] ),
    .X(_0379_));
 sky130_fd_sc_hd__and4_1 _1108_ (.A(\rgb_mixer.debounce2_b.button_hist[0] ),
    .B(\rgb_mixer.debounce2_b.button_hist[1] ),
    .C(\rgb_mixer.debounce2_b.button_hist[2] ),
    .D(\rgb_mixer.debounce2_b.button_hist[3] ),
    .X(_0380_));
 sky130_fd_sc_hd__or4_1 _1109_ (.A(\rgb_mixer.debounce2_b.button_hist[0] ),
    .B(\rgb_mixer.debounce2_b.button_hist[1] ),
    .C(\rgb_mixer.debounce2_b.button_hist[2] ),
    .D(\rgb_mixer.debounce2_b.button_hist[3] ),
    .X(_0381_));
 sky130_fd_sc_hd__or4_1 _1110_ (.A(\rgb_mixer.debounce2_b.button_hist[4] ),
    .B(\rgb_mixer.debounce2_b.button_hist[5] ),
    .C(\rgb_mixer.debounce2_b.button_hist[7] ),
    .D(\rgb_mixer.debounce2_b.button_hist[6] ),
    .X(_0382_));
 sky130_fd_sc_hd__or2_1 _1111_ (.A(_0381_),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__a32o_1 _1112_ (.A1(_0247_),
    .A2(_0379_),
    .A3(_0380_),
    .B1(_0383_),
    .B2(_0024_),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _1113_ (.A(_0269_),
    .B(net4),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _1114_ (.A(_0384_),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _1115_ (.A(\rgb_mixer.debounce2_a.button_hist[0] ),
    .B(_0161_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _1116_ (.A(_0385_),
    .X(_0064_));
 sky130_fd_sc_hd__and2_1 _1117_ (.A(\rgb_mixer.debounce2_a.button_hist[1] ),
    .B(_0370_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _1118_ (.A(_0386_),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _1119_ (.A(\rgb_mixer.debounce2_a.button_hist[2] ),
    .B(_0370_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _1120_ (.A(_0387_),
    .X(_0066_));
 sky130_fd_sc_hd__and2_1 _1121_ (.A(\rgb_mixer.debounce2_a.button_hist[3] ),
    .B(_0370_),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _1122_ (.A(_0388_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_2 _1123_ (.A(_0161_),
    .X(_0389_));
 sky130_fd_sc_hd__and2_1 _1124_ (.A(\rgb_mixer.debounce2_a.button_hist[4] ),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _1125_ (.A(_0390_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _1126_ (.A(\rgb_mixer.debounce2_a.button_hist[5] ),
    .B(_0389_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _1127_ (.A(_0391_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _1128_ (.A(\rgb_mixer.debounce2_a.button_hist[6] ),
    .B(_0389_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _1129_ (.A(_0392_),
    .X(_0070_));
 sky130_fd_sc_hd__and4_1 _1130_ (.A(\rgb_mixer.debounce2_a.button_hist[5] ),
    .B(\rgb_mixer.debounce2_a.button_hist[4] ),
    .C(\rgb_mixer.debounce2_a.button_hist[7] ),
    .D(\rgb_mixer.debounce2_a.button_hist[6] ),
    .X(_0393_));
 sky130_fd_sc_hd__and3_1 _1131_ (.A(\rgb_mixer.debounce2_a.button_hist[1] ),
    .B(\rgb_mixer.debounce2_a.button_hist[2] ),
    .C(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__or3_1 _1132_ (.A(\rgb_mixer.debounce2_a.button_hist[1] ),
    .B(\rgb_mixer.debounce2_a.button_hist[0] ),
    .C(\rgb_mixer.debounce2_a.button_hist[3] ),
    .X(_0395_));
 sky130_fd_sc_hd__or4_1 _1133_ (.A(\rgb_mixer.debounce2_a.button_hist[5] ),
    .B(\rgb_mixer.debounce2_a.button_hist[4] ),
    .C(\rgb_mixer.debounce2_a.button_hist[7] ),
    .D(\rgb_mixer.debounce2_a.button_hist[6] ),
    .X(_0396_));
 sky130_fd_sc_hd__o31a_1 _1134_ (.A1(\rgb_mixer.debounce2_a.button_hist[2] ),
    .A2(_0395_),
    .A3(_0396_),
    .B1(\rgb_mixer.debounce2_a.debounced ),
    .X(_0397_));
 sky130_fd_sc_hd__a32o_1 _1135_ (.A1(\rgb_mixer.debounce2_a.button_hist[3] ),
    .A2(_0064_),
    .A3(_0394_),
    .B1(_0397_),
    .B2(_0247_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _1136_ (.A(_0269_),
    .B(net3),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _1137_ (.A(_0398_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _1138_ (.A(\rgb_mixer.debounce1_b.button_hist[0] ),
    .B(_0160_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _1139_ (.A(_0399_),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _1140_ (.A(\rgb_mixer.debounce1_b.button_hist[1] ),
    .B(_0389_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _1141_ (.A(_0400_),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _1142_ (.A(\rgb_mixer.debounce1_b.button_hist[2] ),
    .B(_0389_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1143_ (.A(_0401_),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _1144_ (.A(\rgb_mixer.debounce1_b.button_hist[3] ),
    .B(_0389_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _1145_ (.A(_0402_),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _1146_ (.A(\rgb_mixer.debounce1_b.button_hist[4] ),
    .B(_0389_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _1147_ (.A(_0403_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _1148_ (.A(\rgb_mixer.debounce1_b.button_hist[5] ),
    .B(_0389_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _1149_ (.A(_0404_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _1150_ (.A(\rgb_mixer.debounce1_b.button_hist[6] ),
    .B(_0389_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _1151_ (.A(_0405_),
    .X(_0079_));
 sky130_fd_sc_hd__and4_1 _1152_ (.A(\rgb_mixer.debounce1_b.button_hist[5] ),
    .B(\rgb_mixer.debounce1_b.button_hist[4] ),
    .C(\rgb_mixer.debounce1_b.button_hist[7] ),
    .D(\rgb_mixer.debounce1_b.button_hist[6] ),
    .X(_0406_));
 sky130_fd_sc_hd__and3_1 _1153_ (.A(\rgb_mixer.debounce1_b.button_hist[1] ),
    .B(\rgb_mixer.debounce1_b.button_hist[2] ),
    .C(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__or3_1 _1154_ (.A(\rgb_mixer.debounce1_b.button_hist[1] ),
    .B(\rgb_mixer.debounce1_b.button_hist[0] ),
    .C(\rgb_mixer.debounce1_b.button_hist[3] ),
    .X(_0408_));
 sky130_fd_sc_hd__or4_1 _1155_ (.A(\rgb_mixer.debounce1_b.button_hist[5] ),
    .B(\rgb_mixer.debounce1_b.button_hist[4] ),
    .C(\rgb_mixer.debounce1_b.button_hist[7] ),
    .D(\rgb_mixer.debounce1_b.button_hist[6] ),
    .X(_0409_));
 sky130_fd_sc_hd__o31a_1 _1156_ (.A1(\rgb_mixer.debounce1_b.button_hist[2] ),
    .A2(_0408_),
    .A3(_0409_),
    .B1(\rgb_mixer.debounce1_b.debounced ),
    .X(_0410_));
 sky130_fd_sc_hd__a32o_1 _1157_ (.A1(\rgb_mixer.debounce1_b.button_hist[3] ),
    .A2(_0073_),
    .A3(_0407_),
    .B1(_0410_),
    .B2(_0247_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _1158_ (.A(_0269_),
    .B(net2),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _1159_ (.A(_0411_),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _1160_ (.A(\rgb_mixer.debounce1_a.button_hist[0] ),
    .B(_0160_),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _1161_ (.A(_0412_),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _1162_ (.A(\rgb_mixer.debounce1_a.button_hist[1] ),
    .B(_0389_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _1163_ (.A(_0413_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_2 _1164_ (.A(_0161_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _1165_ (.A(\rgb_mixer.debounce1_a.button_hist[2] ),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _1166_ (.A(_0415_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _1167_ (.A(\rgb_mixer.debounce1_a.button_hist[3] ),
    .B(_0414_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _1168_ (.A(_0416_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _1169_ (.A(\rgb_mixer.debounce1_a.button_hist[4] ),
    .B(_0414_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _1170_ (.A(_0417_),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _1171_ (.A(\rgb_mixer.debounce1_a.button_hist[5] ),
    .B(_0414_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _1172_ (.A(_0418_),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _1173_ (.A(\rgb_mixer.debounce1_a.button_hist[6] ),
    .B(_0414_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _1174_ (.A(_0419_),
    .X(_0088_));
 sky130_fd_sc_hd__and4_1 _1175_ (.A(\rgb_mixer.debounce1_a.button_hist[5] ),
    .B(\rgb_mixer.debounce1_a.button_hist[4] ),
    .C(\rgb_mixer.debounce1_a.button_hist[7] ),
    .D(\rgb_mixer.debounce1_a.button_hist[6] ),
    .X(_0420_));
 sky130_fd_sc_hd__and3_1 _1176_ (.A(\rgb_mixer.debounce1_a.button_hist[1] ),
    .B(\rgb_mixer.debounce1_a.button_hist[2] ),
    .C(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__or3_1 _1177_ (.A(\rgb_mixer.debounce1_a.button_hist[1] ),
    .B(\rgb_mixer.debounce1_a.button_hist[0] ),
    .C(\rgb_mixer.debounce1_a.button_hist[3] ),
    .X(_0422_));
 sky130_fd_sc_hd__or4_1 _1178_ (.A(\rgb_mixer.debounce1_a.button_hist[5] ),
    .B(\rgb_mixer.debounce1_a.button_hist[4] ),
    .C(\rgb_mixer.debounce1_a.button_hist[7] ),
    .D(\rgb_mixer.debounce1_a.button_hist[6] ),
    .X(_0423_));
 sky130_fd_sc_hd__o31a_1 _1179_ (.A1(\rgb_mixer.debounce1_a.button_hist[2] ),
    .A2(_0422_),
    .A3(_0423_),
    .B1(\rgb_mixer.debounce1_a.debounced ),
    .X(_0424_));
 sky130_fd_sc_hd__a32o_1 _1180_ (.A1(\rgb_mixer.debounce1_a.button_hist[3] ),
    .A2(_0082_),
    .A3(_0421_),
    .B1(_0424_),
    .B2(_0247_),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _1181_ (.A(_0269_),
    .B(net7),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _1182_ (.A(_0425_),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _1183_ (.A(\rgb_mixer.debounce0_b.button_hist[0] ),
    .B(_0160_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _1184_ (.A(_0426_),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _1185_ (.A(\rgb_mixer.debounce0_b.button_hist[1] ),
    .B(_0414_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _1186_ (.A(_0427_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _1187_ (.A(\rgb_mixer.debounce0_b.button_hist[2] ),
    .B(_0414_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _1188_ (.A(_0428_),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _1189_ (.A(\rgb_mixer.debounce0_b.button_hist[3] ),
    .B(_0414_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _1190_ (.A(_0429_),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _1191_ (.A(\rgb_mixer.debounce0_b.button_hist[4] ),
    .B(_0414_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1192_ (.A(_0430_),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _1193_ (.A(\rgb_mixer.debounce0_b.button_hist[5] ),
    .B(_0414_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _1194_ (.A(_0431_),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _1195_ (.A(\rgb_mixer.debounce0_b.button_hist[6] ),
    .B(_0162_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1196_ (.A(_0432_),
    .X(_0097_));
 sky130_fd_sc_hd__and4_1 _1197_ (.A(\rgb_mixer.debounce0_b.button_hist[5] ),
    .B(\rgb_mixer.debounce0_b.button_hist[4] ),
    .C(\rgb_mixer.debounce0_b.button_hist[7] ),
    .D(\rgb_mixer.debounce0_b.button_hist[6] ),
    .X(_0433_));
 sky130_fd_sc_hd__and3_1 _1198_ (.A(\rgb_mixer.debounce0_b.button_hist[1] ),
    .B(\rgb_mixer.debounce0_b.button_hist[2] ),
    .C(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__or3_1 _1199_ (.A(\rgb_mixer.debounce0_b.button_hist[1] ),
    .B(\rgb_mixer.debounce0_b.button_hist[0] ),
    .C(\rgb_mixer.debounce0_b.button_hist[3] ),
    .X(_0435_));
 sky130_fd_sc_hd__or4_1 _1200_ (.A(\rgb_mixer.debounce0_b.button_hist[5] ),
    .B(\rgb_mixer.debounce0_b.button_hist[4] ),
    .C(\rgb_mixer.debounce0_b.button_hist[7] ),
    .D(\rgb_mixer.debounce0_b.button_hist[6] ),
    .X(_0436_));
 sky130_fd_sc_hd__o31a_1 _1201_ (.A1(\rgb_mixer.debounce0_b.button_hist[2] ),
    .A2(_0435_),
    .A3(_0436_),
    .B1(\rgb_mixer.debounce0_b.debounced ),
    .X(_0437_));
 sky130_fd_sc_hd__a32o_1 _1202_ (.A1(\rgb_mixer.debounce0_b.button_hist[3] ),
    .A2(_0091_),
    .A3(_0434_),
    .B1(_0437_),
    .B2(_0247_),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _1203_ (.A(_0269_),
    .B(net6),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _1204_ (.A(_0438_),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _1205_ (.A(\rgb_mixer.debounce0_a.button_hist[0] ),
    .B(_0162_),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _1206_ (.A(_0439_),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _1207_ (.A(\rgb_mixer.debounce0_a.button_hist[1] ),
    .B(_0162_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _1208_ (.A(_0440_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _1209_ (.A(\rgb_mixer.debounce0_a.button_hist[2] ),
    .B(_0162_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _1210_ (.A(_0441_),
    .X(_0102_));
 sky130_fd_sc_hd__and2_1 _1211_ (.A(\rgb_mixer.debounce0_a.button_hist[3] ),
    .B(_0162_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _1212_ (.A(_0442_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _1213_ (.A(\rgb_mixer.debounce0_a.button_hist[4] ),
    .B(_0162_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _1214_ (.A(_0443_),
    .X(_0104_));
 sky130_fd_sc_hd__and2_1 _1215_ (.A(\rgb_mixer.debounce0_a.button_hist[5] ),
    .B(_0162_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _1216_ (.A(_0444_),
    .X(_0105_));
 sky130_fd_sc_hd__and2_1 _1217_ (.A(\rgb_mixer.debounce0_a.button_hist[6] ),
    .B(_0162_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _1218_ (.A(_0445_),
    .X(_0106_));
 sky130_fd_sc_hd__and4_1 _1219_ (.A(\rgb_mixer.debounce0_a.button_hist[5] ),
    .B(\rgb_mixer.debounce0_a.button_hist[4] ),
    .C(\rgb_mixer.debounce0_a.button_hist[7] ),
    .D(\rgb_mixer.debounce0_a.button_hist[6] ),
    .X(_0446_));
 sky130_fd_sc_hd__and4_1 _1220_ (.A(\rgb_mixer.debounce0_a.button_hist[1] ),
    .B(\rgb_mixer.debounce0_a.button_hist[0] ),
    .C(\rgb_mixer.debounce0_a.button_hist[3] ),
    .D(\rgb_mixer.debounce0_a.button_hist[2] ),
    .X(_0447_));
 sky130_fd_sc_hd__or4_1 _1221_ (.A(\rgb_mixer.debounce0_a.button_hist[1] ),
    .B(\rgb_mixer.debounce0_a.button_hist[0] ),
    .C(\rgb_mixer.debounce0_a.button_hist[3] ),
    .D(\rgb_mixer.debounce0_a.button_hist[2] ),
    .X(_0448_));
 sky130_fd_sc_hd__or4_1 _1222_ (.A(\rgb_mixer.debounce0_a.button_hist[5] ),
    .B(\rgb_mixer.debounce0_a.button_hist[4] ),
    .C(\rgb_mixer.debounce0_a.button_hist[7] ),
    .D(\rgb_mixer.debounce0_a.button_hist[6] ),
    .X(_0449_));
 sky130_fd_sc_hd__or2_1 _1223_ (.A(_0448_),
    .B(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__a32o_1 _1224_ (.A1(_0188_),
    .A2(_0446_),
    .A3(_0447_),
    .B1(_0450_),
    .B2(_0061_),
    .X(_0107_));
 sky130_fd_sc_hd__dfxtp_1 _1225_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0000_),
    .Q(\rgb_mixer.pwm2.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1226_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0001_),
    .Q(\rgb_mixer.pwm2.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1227_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0002_),
    .Q(\rgb_mixer.pwm2.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1228_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0003_),
    .Q(\rgb_mixer.pwm2.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1229_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0004_),
    .Q(\rgb_mixer.pwm2.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1230_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0005_),
    .Q(\rgb_mixer.pwm2.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1231_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0006_),
    .Q(\rgb_mixer.pwm2.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1232_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0007_),
    .Q(\rgb_mixer.pwm2.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1233_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0008_),
    .Q(\rgb_mixer.pwm1.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0009_),
    .Q(\rgb_mixer.pwm1.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0010_),
    .Q(\rgb_mixer.pwm1.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1236_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0011_),
    .Q(\rgb_mixer.pwm1.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0012_),
    .Q(\rgb_mixer.pwm1.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1238_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0013_),
    .Q(\rgb_mixer.pwm1.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1239_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0014_),
    .Q(\rgb_mixer.pwm1.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0015_),
    .Q(\rgb_mixer.pwm1.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0016_),
    .Q(\rgb_mixer.pwm0.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0017_),
    .Q(\rgb_mixer.pwm0.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0018_),
    .Q(\rgb_mixer.pwm0.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1244_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0019_),
    .Q(\rgb_mixer.pwm0.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1245_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0020_),
    .Q(\rgb_mixer.pwm0.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0021_),
    .Q(\rgb_mixer.pwm0.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0022_),
    .Q(\rgb_mixer.pwm0.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0023_),
    .Q(\rgb_mixer.pwm0.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0024_),
    .Q(\rgb_mixer.encoder2.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0025_),
    .Q(\rgb_mixer.enc2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0026_),
    .Q(\rgb_mixer.enc2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0027_),
    .Q(\rgb_mixer.enc2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0028_),
    .Q(\rgb_mixer.enc2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0029_),
    .Q(\rgb_mixer.enc2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0030_),
    .Q(\rgb_mixer.enc2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0031_),
    .Q(\rgb_mixer.enc2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1257_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0032_),
    .Q(\rgb_mixer.enc2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0033_),
    .Q(\rgb_mixer.encoder1.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _1259_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0034_),
    .Q(\rgb_mixer.encoder2.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0035_),
    .Q(\rgb_mixer.enc1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0036_),
    .Q(\rgb_mixer.enc1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0037_),
    .Q(\rgb_mixer.enc1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0038_),
    .Q(\rgb_mixer.enc1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0039_),
    .Q(\rgb_mixer.enc1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0040_),
    .Q(\rgb_mixer.enc1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0041_),
    .Q(\rgb_mixer.enc1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0042_),
    .Q(\rgb_mixer.enc1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0043_),
    .Q(\rgb_mixer.encoder0.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0044_),
    .Q(\rgb_mixer.encoder1.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _1270_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0045_),
    .Q(\rgb_mixer.enc0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1271_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0046_),
    .Q(\rgb_mixer.enc0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1272_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0047_),
    .Q(\rgb_mixer.enc0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1273_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0048_),
    .Q(\rgb_mixer.enc0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1274_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0049_),
    .Q(\rgb_mixer.enc0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1275_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0050_),
    .Q(\rgb_mixer.enc0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1276_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0051_),
    .Q(\rgb_mixer.enc0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1277_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0052_),
    .Q(\rgb_mixer.enc0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1278_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0053_),
    .Q(\rgb_mixer.debounce2_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1279_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0054_),
    .Q(\rgb_mixer.debounce2_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1280_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0055_),
    .Q(\rgb_mixer.debounce2_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1281_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0056_),
    .Q(\rgb_mixer.debounce2_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1282_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0057_),
    .Q(\rgb_mixer.debounce2_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1283_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0058_),
    .Q(\rgb_mixer.debounce2_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1284_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0059_),
    .Q(\rgb_mixer.debounce2_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1285_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0060_),
    .Q(\rgb_mixer.debounce2_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1286_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0061_),
    .Q(\rgb_mixer.encoder0.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _1287_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0062_),
    .Q(\rgb_mixer.debounce2_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1288_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0063_),
    .Q(\rgb_mixer.debounce2_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1289_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0064_),
    .Q(\rgb_mixer.debounce2_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1290_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0065_),
    .Q(\rgb_mixer.debounce2_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1291_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0066_),
    .Q(\rgb_mixer.debounce2_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1292_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0067_),
    .Q(\rgb_mixer.debounce2_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1293_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0068_),
    .Q(\rgb_mixer.debounce2_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1294_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0069_),
    .Q(\rgb_mixer.debounce2_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1295_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0070_),
    .Q(\rgb_mixer.debounce2_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1296_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0071_),
    .Q(\rgb_mixer.debounce2_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1297_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0072_),
    .Q(\rgb_mixer.debounce1_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1298_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0073_),
    .Q(\rgb_mixer.debounce1_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1299_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0074_),
    .Q(\rgb_mixer.debounce1_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1300_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0075_),
    .Q(\rgb_mixer.debounce1_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1301_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0076_),
    .Q(\rgb_mixer.debounce1_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1302_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0077_),
    .Q(\rgb_mixer.debounce1_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1303_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0078_),
    .Q(\rgb_mixer.debounce1_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1304_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0079_),
    .Q(\rgb_mixer.debounce1_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1305_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0080_),
    .Q(\rgb_mixer.debounce1_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1306_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0081_),
    .Q(\rgb_mixer.debounce1_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1307_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0082_),
    .Q(\rgb_mixer.debounce1_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1308_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0083_),
    .Q(\rgb_mixer.debounce1_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1309_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0084_),
    .Q(\rgb_mixer.debounce1_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1310_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0085_),
    .Q(\rgb_mixer.debounce1_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1311_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0086_),
    .Q(\rgb_mixer.debounce1_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1312_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0087_),
    .Q(\rgb_mixer.debounce1_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1313_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0088_),
    .Q(\rgb_mixer.debounce1_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1314_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0089_),
    .Q(\rgb_mixer.debounce1_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1315_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0090_),
    .Q(\rgb_mixer.debounce0_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1316_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0091_),
    .Q(\rgb_mixer.debounce0_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1317_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0092_),
    .Q(\rgb_mixer.debounce0_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1318_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0093_),
    .Q(\rgb_mixer.debounce0_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1319_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0094_),
    .Q(\rgb_mixer.debounce0_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1320_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0095_),
    .Q(\rgb_mixer.debounce0_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1321_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0096_),
    .Q(\rgb_mixer.debounce0_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1322_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0097_),
    .Q(\rgb_mixer.debounce0_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1323_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0098_),
    .Q(\rgb_mixer.debounce0_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1324_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0099_),
    .Q(\rgb_mixer.debounce0_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1325_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0100_),
    .Q(\rgb_mixer.debounce0_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1326_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0101_),
    .Q(\rgb_mixer.debounce0_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1327_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0102_),
    .Q(\rgb_mixer.debounce0_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1328_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0103_),
    .Q(\rgb_mixer.debounce0_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1329_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0104_),
    .Q(\rgb_mixer.debounce0_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1330_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0105_),
    .Q(\rgb_mixer.debounce0_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1331_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0106_),
    .Q(\rgb_mixer.debounce0_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1332_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0107_),
    .Q(\rgb_mixer.debounce0_a.debounced ));
 sky130_fd_sc_hd__conb_1 _1438__10 (.LO(net10));
 sky130_fd_sc_hd__conb_1 _1439__11 (.LO(net11));
 sky130_fd_sc_hd__conb_1 _1440__12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 _1441__13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 _1442__14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 _1443__15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 _1444__16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 _1445__17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 _1446__18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 _1447__19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 _1448__20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 _1449__21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 _1450__22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 _1451__23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 _1452__24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 _1453__25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 _1454__26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _1455__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _1456__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _1457__29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _1458__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _1459__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _1460__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _1461__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _1462__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _1463__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _1464__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _1465__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _1466__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _1467__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _1468__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _1469__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _1470__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _1471__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _1472__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _1473__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _1474__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _1475__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _1476__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _1477__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _1478__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _1479__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _1480__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _1481__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _1482__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _1487__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _1488__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _1489__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _1490__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _1491__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _1492__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _1493__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _1494__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _1495__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _1496__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _1497__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _1498__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _1499__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _1500__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _1501__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _1502__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _1503__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _1504__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _1505__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _1506__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _1507__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _1508__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _1509__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _1510__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _1511__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _1512__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _1513__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _1514__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _1515__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _1516__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _1517__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _1518__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _1519__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _1520__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _1521__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _1522__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _1523__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _1524__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _1525__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _1526__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _1527__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _1528__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _1529__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _1530__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _1531__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _1532__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _1533__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _1534__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _1535__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _1536__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _1537__105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 _1538__106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 _1539__107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 _1540__108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 _1541__109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 _1542__110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 _1543__111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 _1544__112 (.LO(net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _1437_ (.A(net9),
    .TE_B(_0451_),
    .Z(la1_data_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1438_ (.A(net10),
    .TE_B(_0452_),
    .Z(la1_data_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1439_ (.A(net11),
    .TE_B(_0453_),
    .Z(la1_data_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1440_ (.A(net12),
    .TE_B(_0454_),
    .Z(la1_data_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1441_ (.A(net13),
    .TE_B(_0455_),
    .Z(la1_data_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1442_ (.A(net14),
    .TE_B(_0456_),
    .Z(la1_data_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1443_ (.A(net15),
    .TE_B(_0457_),
    .Z(la1_data_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1444_ (.A(net16),
    .TE_B(_0458_),
    .Z(la1_data_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1445_ (.A(net17),
    .TE_B(_0459_),
    .Z(la1_data_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1446_ (.A(net18),
    .TE_B(_0460_),
    .Z(la1_data_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1447_ (.A(net19),
    .TE_B(_0461_),
    .Z(la1_data_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1448_ (.A(net20),
    .TE_B(_0462_),
    .Z(la1_data_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1449_ (.A(net21),
    .TE_B(_0463_),
    .Z(la1_data_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1450_ (.A(net22),
    .TE_B(_0464_),
    .Z(la1_data_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1451_ (.A(net23),
    .TE_B(_0465_),
    .Z(la1_data_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1452_ (.A(net24),
    .TE_B(_0466_),
    .Z(la1_data_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1453_ (.A(net25),
    .TE_B(_0467_),
    .Z(la1_data_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1454_ (.A(net26),
    .TE_B(_0468_),
    .Z(la1_data_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1455_ (.A(net27),
    .TE_B(_0469_),
    .Z(la1_data_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1456_ (.A(net28),
    .TE_B(_0470_),
    .Z(la1_data_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1457_ (.A(net29),
    .TE_B(_0471_),
    .Z(la1_data_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1458_ (.A(net30),
    .TE_B(_0472_),
    .Z(la1_data_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1459_ (.A(net31),
    .TE_B(_0473_),
    .Z(la1_data_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1460_ (.A(net32),
    .TE_B(_0474_),
    .Z(la1_data_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1461_ (.A(net33),
    .TE_B(_0475_),
    .Z(la1_data_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1462_ (.A(net34),
    .TE_B(_0476_),
    .Z(la1_data_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1463_ (.A(net35),
    .TE_B(_0477_),
    .Z(la1_data_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1464_ (.A(net36),
    .TE_B(_0478_),
    .Z(la1_data_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1465_ (.A(net37),
    .TE_B(_0479_),
    .Z(la1_data_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1466_ (.A(net38),
    .TE_B(_0480_),
    .Z(la1_data_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1467_ (.A(net39),
    .TE_B(_0481_),
    .Z(la1_data_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1468_ (.A(net40),
    .TE_B(_0482_),
    .Z(la1_data_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1469_ (.A(net41),
    .TE_B(_0483_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1470_ (.A(net42),
    .TE_B(_0484_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1471_ (.A(net43),
    .TE_B(_0485_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1472_ (.A(net44),
    .TE_B(_0486_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1473_ (.A(net45),
    .TE_B(_0487_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1474_ (.A(net46),
    .TE_B(_0488_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1475_ (.A(net47),
    .TE_B(_0489_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1476_ (.A(net48),
    .TE_B(_0490_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1477_ (.A(net49),
    .TE_B(_0491_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1478_ (.A(net50),
    .TE_B(_0492_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1479_ (.A(net51),
    .TE_B(_0493_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1480_ (.A(net52),
    .TE_B(_0494_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1481_ (.A(net53),
    .TE_B(_0495_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1482_ (.A(net54),
    .TE_B(_0496_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1483_ (.A(\rgb_mixer.pwm0.out ),
    .TE_B(_0497_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1484_ (.A(\rgb_mixer.pwm1.out ),
    .TE_B(_0498_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1485_ (.A(\rgb_mixer.pwm2.out ),
    .TE_B(_0499_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1486_ (.A(net8),
    .TE_B(_0500_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1487_ (.A(net55),
    .TE_B(_0501_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1488_ (.A(net56),
    .TE_B(_0502_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1489_ (.A(net57),
    .TE_B(_0503_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1490_ (.A(net58),
    .TE_B(_0504_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1491_ (.A(net59),
    .TE_B(_0505_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1492_ (.A(net60),
    .TE_B(_0506_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1493_ (.A(net61),
    .TE_B(_0507_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1494_ (.A(net62),
    .TE_B(_0508_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1495_ (.A(net63),
    .TE_B(_0509_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1496_ (.A(net64),
    .TE_B(_0510_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1497_ (.A(net65),
    .TE_B(_0511_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1498_ (.A(net66),
    .TE_B(_0512_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1499_ (.A(net67),
    .TE_B(_0513_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1500_ (.A(net68),
    .TE_B(_0514_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1501_ (.A(net69),
    .TE_B(_0515_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _1502_ (.A(net70),
    .TE_B(_0516_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _1503_ (.A(net71),
    .TE_B(_0517_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _1504_ (.A(net72),
    .TE_B(_0518_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _1505_ (.A(net73),
    .TE_B(_0519_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _1506_ (.A(net74),
    .TE_B(_0520_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _1507_ (.A(net75),
    .TE_B(_0521_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _1508_ (.A(net76),
    .TE_B(_0522_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _1509_ (.A(net77),
    .TE_B(_0523_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _1510_ (.A(net78),
    .TE_B(_0524_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _1511_ (.A(net79),
    .TE_B(_0525_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _1512_ (.A(net80),
    .TE_B(_0526_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _1513_ (.A(net81),
    .TE_B(_0527_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _1514_ (.A(net82),
    .TE_B(_0528_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _1515_ (.A(net83),
    .TE_B(_0529_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _1516_ (.A(net84),
    .TE_B(_0530_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _1517_ (.A(net85),
    .TE_B(_0531_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _1518_ (.A(net86),
    .TE_B(_0532_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _1519_ (.A(net87),
    .TE_B(_0533_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _1520_ (.A(net88),
    .TE_B(_0534_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _1521_ (.A(net89),
    .TE_B(_0535_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _1522_ (.A(net90),
    .TE_B(_0536_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _1523_ (.A(net91),
    .TE_B(_0537_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _1524_ (.A(net92),
    .TE_B(_0538_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _1525_ (.A(net93),
    .TE_B(_0539_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _1526_ (.A(net94),
    .TE_B(_0540_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _1527_ (.A(net95),
    .TE_B(_0541_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _1528_ (.A(net96),
    .TE_B(_0542_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _1529_ (.A(net97),
    .TE_B(_0543_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _1530_ (.A(net98),
    .TE_B(_0544_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _1531_ (.A(net99),
    .TE_B(_0545_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _1532_ (.A(net100),
    .TE_B(_0546_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _1533_ (.A(net101),
    .TE_B(_0547_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _1534_ (.A(net102),
    .TE_B(_0548_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _1535_ (.A(net103),
    .TE_B(_0549_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _1536_ (.A(net104),
    .TE_B(_0550_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _1537_ (.A(net105),
    .TE_B(_0551_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _1538_ (.A(net106),
    .TE_B(_0552_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _1539_ (.A(net107),
    .TE_B(_0553_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _1540_ (.A(net108),
    .TE_B(_0554_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _1541_ (.A(net109),
    .TE_B(_0555_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _1542_ (.A(net110),
    .TE_B(_0556_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _1543_ (.A(net111),
    .TE_B(_0557_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _1544_ (.A(net112),
    .TE_B(_0558_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(io_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[8]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[9]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(la1_data_in[0]),
    .X(net8));
 sky130_fd_sc_hd__conb_1 _1437__9 (.LO(net9));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net7));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_510 ();
endmodule

