magic
tech sky130A
magscale 1 2
timestamp 1672827330
<< viali >>
rect 47225 47073 47259 47107
rect 1961 47005 1995 47039
rect 2697 47005 2731 47039
rect 4537 47005 4571 47039
rect 5181 47005 5215 47039
rect 5641 47005 5675 47039
rect 6745 47005 6779 47039
rect 7389 47005 7423 47039
rect 8033 47005 8067 47039
rect 9321 47005 9355 47039
rect 12541 47005 12575 47039
rect 14565 47005 14599 47039
rect 15209 47005 15243 47039
rect 23029 47005 23063 47039
rect 25329 47005 25363 47039
rect 27353 47005 27387 47039
rect 27997 47005 28031 47039
rect 29101 47005 29135 47039
rect 29929 47005 29963 47039
rect 33241 47005 33275 47039
rect 38301 47005 38335 47039
rect 41613 47005 41647 47039
rect 44649 47005 44683 47039
rect 45385 47005 45419 47039
rect 47777 47005 47811 47039
rect 3249 46937 3283 46971
rect 45569 46937 45603 46971
rect 47869 46937 47903 46971
rect 2053 46869 2087 46903
rect 5733 46869 5767 46903
rect 7849 46869 7883 46903
rect 9137 46869 9171 46903
rect 27813 46869 27847 46903
rect 2053 46597 2087 46631
rect 6745 46597 6779 46631
rect 47225 46597 47259 46631
rect 1869 46529 1903 46563
rect 4169 46529 4203 46563
rect 6561 46529 6595 46563
rect 12173 46529 12207 46563
rect 14473 46529 14507 46563
rect 22477 46529 22511 46563
rect 24777 46529 24811 46563
rect 27169 46529 27203 46563
rect 29469 46529 29503 46563
rect 32965 46529 32999 46563
rect 39773 46529 39807 46563
rect 42625 46529 42659 46563
rect 45385 46529 45419 46563
rect 2789 46461 2823 46495
rect 4353 46461 4387 46495
rect 4721 46461 4755 46495
rect 7021 46461 7055 46495
rect 12357 46461 12391 46495
rect 12909 46461 12943 46495
rect 14657 46461 14691 46495
rect 15485 46461 15519 46495
rect 22661 46461 22695 46495
rect 23213 46461 23247 46495
rect 24961 46461 24995 46495
rect 25789 46461 25823 46495
rect 27353 46461 27387 46495
rect 27629 46461 27663 46495
rect 29653 46461 29687 46495
rect 29929 46461 29963 46495
rect 33149 46461 33183 46495
rect 33517 46461 33551 46495
rect 36553 46461 36587 46495
rect 37473 46461 37507 46495
rect 37657 46461 37691 46495
rect 37933 46461 37967 46495
rect 39957 46461 39991 46495
rect 40233 46461 40267 46495
rect 42809 46461 42843 46495
rect 43085 46461 43119 46495
rect 45569 46461 45603 46495
rect 10701 46325 10735 46359
rect 35817 46325 35851 46359
rect 47961 46325 47995 46359
rect 22937 46121 22971 46155
rect 26985 46121 27019 46155
rect 29101 46121 29135 46155
rect 33241 46121 33275 46155
rect 38025 46121 38059 46155
rect 44557 46121 44591 46155
rect 48145 46121 48179 46155
rect 16681 46053 16715 46087
rect 44005 46053 44039 46087
rect 1777 45985 1811 46019
rect 2789 45985 2823 46019
rect 4905 45985 4939 46019
rect 5641 45985 5675 46019
rect 6101 45985 6135 46019
rect 10425 45985 10459 46019
rect 11069 45985 11103 46019
rect 14289 45985 14323 46019
rect 14841 45985 14875 46019
rect 25145 45985 25179 46019
rect 29745 45985 29779 46019
rect 30389 45985 30423 46019
rect 35541 45985 35575 46019
rect 36093 45985 36127 46019
rect 40601 45985 40635 46019
rect 45753 45985 45787 46019
rect 47133 45985 47167 46019
rect 1593 45917 1627 45951
rect 4353 45917 4387 45951
rect 13093 45917 13127 45951
rect 13553 45917 13587 45951
rect 16589 45917 16623 45951
rect 22845 45917 22879 45951
rect 24041 45917 24075 45951
rect 24593 45917 24627 45951
rect 26893 45917 26927 45951
rect 29009 45917 29043 45951
rect 33149 45917 33183 45951
rect 37933 45917 37967 45951
rect 40141 45917 40175 45951
rect 44465 45917 44499 45951
rect 48053 45917 48087 45951
rect 5825 45849 5859 45883
rect 10609 45849 10643 45883
rect 13645 45849 13679 45883
rect 14473 45849 14507 45883
rect 24777 45849 24811 45883
rect 29929 45849 29963 45883
rect 35725 45849 35759 45883
rect 40325 45849 40359 45883
rect 45937 45849 45971 45883
rect 6653 45577 6687 45611
rect 10609 45577 10643 45611
rect 24501 45577 24535 45611
rect 25329 45577 25363 45611
rect 29837 45577 29871 45611
rect 35725 45577 35759 45611
rect 12449 45509 12483 45543
rect 13093 45509 13127 45543
rect 13829 45509 13863 45543
rect 36645 45509 36679 45543
rect 41613 45509 41647 45543
rect 45569 45509 45603 45543
rect 4721 45441 4755 45475
rect 6561 45441 6595 45475
rect 10517 45441 10551 45475
rect 12357 45441 12391 45475
rect 13001 45441 13035 45475
rect 13645 45441 13679 45475
rect 24409 45441 24443 45475
rect 25237 45441 25271 45475
rect 29745 45441 29779 45475
rect 35633 45441 35667 45475
rect 36553 45441 36587 45475
rect 40417 45441 40451 45475
rect 41521 45441 41555 45475
rect 2237 45373 2271 45407
rect 2421 45373 2455 45407
rect 2973 45373 3007 45407
rect 4997 45373 5031 45407
rect 14197 45373 14231 45407
rect 44925 45373 44959 45407
rect 45385 45373 45419 45407
rect 46857 45373 46891 45407
rect 1777 45237 1811 45271
rect 47961 45237 47995 45271
rect 4445 45033 4479 45067
rect 40325 45033 40359 45067
rect 45845 45033 45879 45067
rect 46489 44897 46523 44931
rect 48237 44897 48271 44931
rect 1777 44829 1811 44863
rect 2605 44829 2639 44863
rect 4353 44829 4387 44863
rect 4997 44829 5031 44863
rect 40233 44829 40267 44863
rect 45753 44829 45787 44863
rect 3249 44761 3283 44795
rect 5825 44761 5859 44795
rect 46673 44761 46707 44795
rect 1869 44693 1903 44727
rect 1685 44489 1719 44523
rect 46489 44489 46523 44523
rect 2421 44421 2455 44455
rect 7389 44421 7423 44455
rect 1593 44353 1627 44387
rect 2237 44353 2271 44387
rect 4537 44353 4571 44387
rect 6561 44353 6595 44387
rect 46397 44353 46431 44387
rect 48329 44353 48363 44387
rect 2789 44285 2823 44319
rect 5457 44285 5491 44319
rect 47225 44149 47259 44183
rect 48145 44149 48179 44183
rect 4077 43945 4111 43979
rect 2789 43809 2823 43843
rect 5549 43809 5583 43843
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 1593 43741 1627 43775
rect 3985 43741 4019 43775
rect 5089 43741 5123 43775
rect 27077 43741 27111 43775
rect 27169 43741 27203 43775
rect 1777 43673 1811 43707
rect 46673 43673 46707 43707
rect 27353 43605 27387 43639
rect 2605 43401 2639 43435
rect 47133 43401 47167 43435
rect 22293 43333 22327 43367
rect 2053 43265 2087 43299
rect 2513 43265 2547 43299
rect 3893 43265 3927 43299
rect 22845 43265 22879 43299
rect 23673 43265 23707 43299
rect 24133 43265 24167 43299
rect 27353 43265 27387 43299
rect 28457 43265 28491 43299
rect 28724 43265 28758 43299
rect 30481 43265 30515 43299
rect 35909 43265 35943 43299
rect 47041 43265 47075 43299
rect 47777 43265 47811 43299
rect 4629 43197 4663 43231
rect 22661 43197 22695 43231
rect 23857 43197 23891 43231
rect 23029 43129 23063 43163
rect 23489 43061 23523 43095
rect 27169 43061 27203 43095
rect 29837 43061 29871 43095
rect 30297 43061 30331 43095
rect 35725 43061 35759 43095
rect 47869 43061 47903 43095
rect 2421 42721 2455 42755
rect 3065 42721 3099 42755
rect 4721 42721 4755 42755
rect 29745 42721 29779 42755
rect 46673 42721 46707 42755
rect 48237 42721 48271 42755
rect 1777 42653 1811 42687
rect 4445 42653 4479 42687
rect 23673 42653 23707 42687
rect 27537 42653 27571 42687
rect 28457 42653 28491 42687
rect 28641 42653 28675 42687
rect 30012 42653 30046 42687
rect 31585 42653 31619 42687
rect 35081 42653 35115 42687
rect 35817 42653 35851 42687
rect 36073 42653 36107 42687
rect 46029 42653 46063 42687
rect 46489 42653 46523 42687
rect 31852 42585 31886 42619
rect 1593 42517 1627 42551
rect 23489 42517 23523 42551
rect 27353 42517 27387 42551
rect 28825 42517 28859 42551
rect 31125 42517 31159 42551
rect 32965 42517 32999 42551
rect 34897 42517 34931 42551
rect 37197 42517 37231 42551
rect 32965 42313 32999 42347
rect 36093 42313 36127 42347
rect 24470 42245 24504 42279
rect 30113 42245 30147 42279
rect 37841 42245 37875 42279
rect 23581 42177 23615 42211
rect 24225 42177 24259 42211
rect 27169 42177 27203 42211
rect 27425 42177 27459 42211
rect 29193 42177 29227 42211
rect 29837 42177 29871 42211
rect 29929 42177 29963 42211
rect 31125 42177 31159 42211
rect 31217 42177 31251 42211
rect 32505 42177 32539 42211
rect 33149 42177 33183 42211
rect 33885 42177 33919 42211
rect 34152 42177 34186 42211
rect 35909 42177 35943 42211
rect 36921 42177 36955 42211
rect 37657 42177 37691 42211
rect 38485 42177 38519 42211
rect 40049 42177 40083 42211
rect 42892 42177 42926 42211
rect 47777 42177 47811 42211
rect 31401 42109 31435 42143
rect 35725 42109 35759 42143
rect 37473 42109 37507 42143
rect 39865 42109 39899 42143
rect 42625 42109 42659 42143
rect 29009 42041 29043 42075
rect 23397 41973 23431 42007
rect 25605 41973 25639 42007
rect 28549 41973 28583 42007
rect 32321 41973 32355 42007
rect 35265 41973 35299 42007
rect 36737 41973 36771 42007
rect 38301 41973 38335 42007
rect 40233 41973 40267 42007
rect 44005 41973 44039 42007
rect 47225 41973 47259 42007
rect 47869 41973 47903 42007
rect 25973 41769 26007 41803
rect 28089 41769 28123 41803
rect 28917 41769 28951 41803
rect 35265 41769 35299 41803
rect 38577 41769 38611 41803
rect 43545 41769 43579 41803
rect 30573 41701 30607 41735
rect 38209 41633 38243 41667
rect 46489 41633 46523 41667
rect 46673 41633 46707 41667
rect 48237 41633 48271 41667
rect 2329 41565 2363 41599
rect 24593 41565 24627 41599
rect 26709 41565 26743 41599
rect 28641 41565 28675 41599
rect 28733 41565 28767 41599
rect 30757 41565 30791 41599
rect 31585 41565 31619 41599
rect 34897 41565 34931 41599
rect 35081 41565 35115 41599
rect 36369 41565 36403 41599
rect 38393 41565 38427 41599
rect 42717 41565 42751 41599
rect 42901 41565 42935 41599
rect 43085 41565 43119 41599
rect 43729 41565 43763 41599
rect 45385 41565 45419 41599
rect 24838 41497 24872 41531
rect 26976 41497 27010 41531
rect 30849 41497 30883 41531
rect 31125 41497 31159 41531
rect 31852 41497 31886 41531
rect 36636 41497 36670 41531
rect 30941 41429 30975 41463
rect 32965 41429 32999 41463
rect 37749 41429 37783 41463
rect 45201 41429 45235 41463
rect 32689 41225 32723 41259
rect 30573 41157 30607 41191
rect 38454 41157 38488 41191
rect 44916 41157 44950 41191
rect 2053 41089 2087 41123
rect 24225 41089 24259 41123
rect 24492 41089 24526 41123
rect 30849 41089 30883 41123
rect 32413 41089 32447 41123
rect 32505 41089 32539 41123
rect 33977 41089 34011 41123
rect 36461 41089 36495 41123
rect 36737 41089 36771 41123
rect 40233 41089 40267 41123
rect 41245 41089 41279 41123
rect 41889 41089 41923 41123
rect 42809 41089 42843 41123
rect 43085 41089 43119 41123
rect 44649 41089 44683 41123
rect 47777 41089 47811 41123
rect 2237 41021 2271 41055
rect 2789 41021 2823 41055
rect 30665 41021 30699 41055
rect 36553 41021 36587 41055
rect 38209 41021 38243 41055
rect 41705 41021 41739 41055
rect 42901 41021 42935 41055
rect 39589 40953 39623 40987
rect 25605 40885 25639 40919
rect 30573 40885 30607 40919
rect 31033 40885 31067 40919
rect 33793 40885 33827 40919
rect 36553 40885 36587 40919
rect 36921 40885 36955 40919
rect 40049 40885 40083 40919
rect 41061 40885 41095 40919
rect 42073 40885 42107 40919
rect 43085 40885 43119 40919
rect 43269 40885 43303 40919
rect 46029 40885 46063 40919
rect 47225 40885 47259 40919
rect 47869 40885 47903 40919
rect 2421 40681 2455 40715
rect 23857 40681 23891 40715
rect 28549 40681 28583 40715
rect 29929 40681 29963 40715
rect 34345 40681 34379 40715
rect 35725 40681 35759 40715
rect 42257 40681 42291 40715
rect 45569 40681 45603 40715
rect 36921 40613 36955 40647
rect 24961 40545 24995 40579
rect 32965 40545 32999 40579
rect 40877 40545 40911 40579
rect 46489 40545 46523 40579
rect 46673 40545 46707 40579
rect 48237 40545 48271 40579
rect 2329 40477 2363 40511
rect 24041 40477 24075 40511
rect 24685 40477 24719 40511
rect 24777 40477 24811 40511
rect 28549 40477 28583 40511
rect 28733 40477 28767 40511
rect 33232 40477 33266 40511
rect 37473 40477 37507 40511
rect 39405 40477 39439 40511
rect 40049 40477 40083 40511
rect 40233 40477 40267 40511
rect 41144 40477 41178 40511
rect 42717 40477 42751 40511
rect 45293 40477 45327 40511
rect 45385 40477 45419 40511
rect 29745 40409 29779 40443
rect 29961 40409 29995 40443
rect 35541 40409 35575 40443
rect 35757 40409 35791 40443
rect 37105 40409 37139 40443
rect 37289 40409 37323 40443
rect 40417 40409 40451 40443
rect 42984 40409 43018 40443
rect 28917 40341 28951 40375
rect 30113 40341 30147 40375
rect 35909 40341 35943 40375
rect 37197 40341 37231 40375
rect 39221 40341 39255 40375
rect 44097 40341 44131 40375
rect 25053 40137 25087 40171
rect 27997 40137 28031 40171
rect 30021 40137 30055 40171
rect 34529 40137 34563 40171
rect 40049 40137 40083 40171
rect 42901 40137 42935 40171
rect 46121 40137 46155 40171
rect 28886 40069 28920 40103
rect 35541 40069 35575 40103
rect 35679 40069 35713 40103
rect 36277 40069 36311 40103
rect 38936 40069 38970 40103
rect 42993 40069 43027 40103
rect 23940 40001 23974 40035
rect 25605 40001 25639 40035
rect 25789 40001 25823 40035
rect 28181 40001 28215 40035
rect 30665 40001 30699 40035
rect 30849 40001 30883 40035
rect 30941 40001 30975 40035
rect 33149 40001 33183 40035
rect 33416 40001 33450 40035
rect 35358 40023 35392 40057
rect 35449 40001 35483 40035
rect 36461 40001 36495 40035
rect 36645 40001 36679 40035
rect 36737 40001 36771 40035
rect 41613 40001 41647 40035
rect 41797 40001 41831 40035
rect 42809 40001 42843 40035
rect 44097 40001 44131 40035
rect 45008 40001 45042 40035
rect 47777 40001 47811 40035
rect 23673 39933 23707 39967
rect 28641 39933 28675 39967
rect 30757 39933 30791 39967
rect 35817 39933 35851 39967
rect 38669 39933 38703 39967
rect 41429 39933 41463 39967
rect 42625 39933 42659 39967
rect 43913 39933 43947 39967
rect 44741 39933 44775 39967
rect 36553 39865 36587 39899
rect 25973 39797 26007 39831
rect 30481 39797 30515 39831
rect 35173 39797 35207 39831
rect 43177 39797 43211 39831
rect 44281 39797 44315 39831
rect 47225 39797 47259 39831
rect 47869 39797 47903 39831
rect 23857 39593 23891 39627
rect 30113 39593 30147 39627
rect 32873 39593 32907 39627
rect 34253 39593 34287 39627
rect 35081 39593 35115 39627
rect 35449 39593 35483 39627
rect 42349 39593 42383 39627
rect 45201 39593 45235 39627
rect 24961 39457 24995 39491
rect 27445 39457 27479 39491
rect 46489 39457 46523 39491
rect 46673 39457 46707 39491
rect 48145 39457 48179 39491
rect 24041 39389 24075 39423
rect 24685 39389 24719 39423
rect 24777 39389 24811 39423
rect 25513 39389 25547 39423
rect 27629 39389 27663 39423
rect 28457 39389 28491 39423
rect 28641 39389 28675 39423
rect 28917 39389 28951 39423
rect 29745 39389 29779 39423
rect 29929 39389 29963 39423
rect 31953 39389 31987 39423
rect 32137 39389 32171 39423
rect 32321 39389 32355 39423
rect 33057 39389 33091 39423
rect 33977 39389 34011 39423
rect 34069 39389 34103 39423
rect 35081 39389 35115 39423
rect 35173 39389 35207 39423
rect 38117 39389 38151 39423
rect 38384 39389 38418 39423
rect 42533 39389 42567 39423
rect 45385 39389 45419 39423
rect 25780 39321 25814 39355
rect 28549 39321 28583 39355
rect 28779 39321 28813 39355
rect 36737 39321 36771 39355
rect 26893 39253 26927 39287
rect 27813 39253 27847 39287
rect 28273 39253 28307 39287
rect 36829 39253 36863 39287
rect 39497 39253 39531 39287
rect 25697 39049 25731 39083
rect 25789 39049 25823 39083
rect 26433 39049 26467 39083
rect 29469 39049 29503 39083
rect 32505 39049 32539 39083
rect 36829 39049 36863 39083
rect 39313 39049 39347 39083
rect 44649 39049 44683 39083
rect 45201 39049 45235 39083
rect 25421 38981 25455 39015
rect 25605 38981 25639 39015
rect 28356 38981 28390 39015
rect 35716 38981 35750 39015
rect 43361 38981 43395 39015
rect 43545 38981 43579 39015
rect 46090 38981 46124 39015
rect 26617 38913 26651 38947
rect 28089 38913 28123 38947
rect 31217 38913 31251 38947
rect 32321 38913 32355 38947
rect 33149 38913 33183 38947
rect 37749 38913 37783 38947
rect 39221 38913 39255 38947
rect 44189 38913 44223 38947
rect 44465 38913 44499 38947
rect 45385 38913 45419 38947
rect 35449 38845 35483 38879
rect 37933 38845 37967 38879
rect 44373 38845 44407 38879
rect 45845 38845 45879 38879
rect 25973 38709 26007 38743
rect 31033 38709 31067 38743
rect 33241 38709 33275 38743
rect 43729 38709 43763 38743
rect 44281 38709 44315 38743
rect 47225 38709 47259 38743
rect 47961 38709 47995 38743
rect 25605 38505 25639 38539
rect 28549 38505 28583 38539
rect 40049 38505 40083 38539
rect 45569 38505 45603 38539
rect 32229 38437 32263 38471
rect 44097 38437 44131 38471
rect 25697 38369 25731 38403
rect 30849 38369 30883 38403
rect 32689 38369 32723 38403
rect 36921 38369 36955 38403
rect 48053 38369 48087 38403
rect 24777 38301 24811 38335
rect 25789 38301 25823 38335
rect 28733 38301 28767 38335
rect 31116 38301 31150 38335
rect 32873 38301 32907 38335
rect 33057 38301 33091 38335
rect 33701 38301 33735 38335
rect 37105 38301 37139 38335
rect 38945 38301 38979 38335
rect 39037 38301 39071 38335
rect 39221 38301 39255 38335
rect 40233 38301 40267 38335
rect 40693 38301 40727 38335
rect 42717 38301 42751 38335
rect 42809 38301 42843 38335
rect 43177 38301 43211 38335
rect 44281 38301 44315 38335
rect 44373 38301 44407 38335
rect 45201 38301 45235 38335
rect 45385 38301 45419 38335
rect 46489 38301 46523 38335
rect 25513 38233 25547 38267
rect 40960 38233 40994 38267
rect 42533 38233 42567 38267
rect 42901 38233 42935 38267
rect 43039 38233 43073 38267
rect 44649 38233 44683 38267
rect 46673 38233 46707 38267
rect 24593 38165 24627 38199
rect 25973 38165 26007 38199
rect 33517 38165 33551 38199
rect 37289 38165 37323 38199
rect 42073 38165 42107 38199
rect 44465 38165 44499 38199
rect 24961 37961 24995 37995
rect 29469 37961 29503 37995
rect 31401 37961 31435 37995
rect 36737 37961 36771 37995
rect 43085 37961 43119 37995
rect 45109 37961 45143 37995
rect 46121 37961 46155 37995
rect 46857 37961 46891 37995
rect 23848 37893 23882 37927
rect 32864 37893 32898 37927
rect 39948 37893 39982 37927
rect 43974 37893 44008 37927
rect 28089 37825 28123 37859
rect 28356 37825 28390 37859
rect 31217 37825 31251 37859
rect 32597 37825 32631 37859
rect 36921 37825 36955 37859
rect 37729 37825 37763 37859
rect 39681 37825 39715 37859
rect 43269 37825 43303 37859
rect 46305 37825 46339 37859
rect 46765 37825 46799 37859
rect 47777 37825 47811 37859
rect 23581 37757 23615 37791
rect 31033 37757 31067 37791
rect 37473 37757 37507 37791
rect 43729 37757 43763 37791
rect 33977 37621 34011 37655
rect 38853 37621 38887 37655
rect 41061 37621 41095 37655
rect 47869 37621 47903 37655
rect 24041 37417 24075 37451
rect 31677 37417 31711 37451
rect 36185 37417 36219 37451
rect 37933 37417 37967 37451
rect 45661 37417 45695 37451
rect 45845 37417 45879 37451
rect 26249 37349 26283 37383
rect 33057 37349 33091 37383
rect 43453 37349 43487 37383
rect 23673 37281 23707 37315
rect 24593 37281 24627 37315
rect 26157 37281 26191 37315
rect 27997 37281 28031 37315
rect 33609 37281 33643 37315
rect 35541 37281 35575 37315
rect 40417 37281 40451 37315
rect 43913 37281 43947 37315
rect 48237 37281 48271 37315
rect 23857 37213 23891 37247
rect 24777 37213 24811 37247
rect 26065 37213 26099 37247
rect 26341 37213 26375 37247
rect 28181 37213 28215 37247
rect 30297 37213 30331 37247
rect 32321 37213 32355 37247
rect 33333 37213 33367 37247
rect 35081 37213 35115 37247
rect 36001 37213 36035 37247
rect 36093 37213 36127 37247
rect 40049 37213 40083 37247
rect 40325 37213 40359 37247
rect 41153 37213 41187 37247
rect 42073 37213 42107 37247
rect 44097 37213 44131 37247
rect 44281 37213 44315 37247
rect 46489 37213 46523 37247
rect 30564 37145 30598 37179
rect 33425 37145 33459 37179
rect 35173 37145 35207 37179
rect 35265 37145 35299 37179
rect 35403 37145 35437 37179
rect 37841 37145 37875 37179
rect 40534 37145 40568 37179
rect 41429 37145 41463 37179
rect 42340 37145 42374 37179
rect 45477 37145 45511 37179
rect 46673 37145 46707 37179
rect 24961 37077 24995 37111
rect 25881 37077 25915 37111
rect 28365 37077 28399 37111
rect 32137 37077 32171 37111
rect 33241 37077 33275 37111
rect 34897 37077 34931 37111
rect 36369 37077 36403 37111
rect 40693 37077 40727 37111
rect 45687 37077 45721 37111
rect 25171 36873 25205 36907
rect 30481 36873 30515 36907
rect 31769 36873 31803 36907
rect 35725 36873 35759 36907
rect 36185 36873 36219 36907
rect 40325 36873 40359 36907
rect 42625 36873 42659 36907
rect 24961 36805 24995 36839
rect 26157 36805 26191 36839
rect 26275 36805 26309 36839
rect 34612 36805 34646 36839
rect 39037 36805 39071 36839
rect 24317 36737 24351 36771
rect 25973 36737 26007 36771
rect 26065 36737 26099 36771
rect 27436 36737 27470 36771
rect 30389 36737 30423 36771
rect 31585 36737 31619 36771
rect 33149 36737 33183 36771
rect 33333 36737 33367 36771
rect 33425 36737 33459 36771
rect 34345 36737 34379 36771
rect 36369 36737 36403 36771
rect 36461 36737 36495 36771
rect 36645 36737 36679 36771
rect 37657 36737 37691 36771
rect 41429 36737 41463 36771
rect 42809 36737 42843 36771
rect 47777 36737 47811 36771
rect 24133 36669 24167 36703
rect 26433 36669 26467 36703
rect 27169 36669 27203 36703
rect 31401 36669 31435 36703
rect 37473 36669 37507 36703
rect 41245 36669 41279 36703
rect 25329 36601 25363 36635
rect 36553 36601 36587 36635
rect 24501 36533 24535 36567
rect 25145 36533 25179 36567
rect 25789 36533 25823 36567
rect 28549 36533 28583 36567
rect 33425 36533 33459 36567
rect 33609 36533 33643 36567
rect 37841 36533 37875 36567
rect 41613 36533 41647 36567
rect 47225 36533 47259 36567
rect 47869 36533 47903 36567
rect 28273 36329 28307 36363
rect 32505 36329 32539 36363
rect 39129 36261 39163 36295
rect 40325 36261 40359 36295
rect 38853 36193 38887 36227
rect 46489 36193 46523 36227
rect 46673 36193 46707 36227
rect 48237 36193 48271 36227
rect 23397 36125 23431 36159
rect 24041 36125 24075 36159
rect 28457 36125 28491 36159
rect 35449 36125 35483 36159
rect 40049 36125 40083 36159
rect 40969 36125 41003 36159
rect 41153 36125 41187 36159
rect 41613 36125 41647 36159
rect 44097 36125 44131 36159
rect 44281 36125 44315 36159
rect 26065 36057 26099 36091
rect 31217 36057 31251 36091
rect 35716 36057 35750 36091
rect 43361 36057 43395 36091
rect 23213 35989 23247 36023
rect 23857 35989 23891 36023
rect 27353 35989 27387 36023
rect 36829 35989 36863 36023
rect 39313 35989 39347 36023
rect 40509 35989 40543 36023
rect 41061 35989 41095 36023
rect 44189 35989 44223 36023
rect 25973 35785 26007 35819
rect 27537 35785 27571 35819
rect 33701 35785 33735 35819
rect 34729 35785 34763 35819
rect 34897 35785 34931 35819
rect 35909 35785 35943 35819
rect 41889 35785 41923 35819
rect 45017 35785 45051 35819
rect 24838 35717 24872 35751
rect 34529 35717 34563 35751
rect 46857 35717 46891 35751
rect 27169 35649 27203 35683
rect 27353 35649 27387 35683
rect 29193 35649 29227 35683
rect 29449 35649 29483 35683
rect 32321 35649 32355 35683
rect 32588 35649 32622 35683
rect 36093 35649 36127 35683
rect 38485 35649 38519 35683
rect 38577 35649 38611 35683
rect 38853 35649 38887 35683
rect 39313 35649 39347 35683
rect 39497 35649 39531 35683
rect 39589 35649 39623 35683
rect 39865 35649 39899 35683
rect 40693 35649 40727 35683
rect 40785 35649 40819 35683
rect 40969 35649 41003 35683
rect 41061 35649 41095 35683
rect 41521 35649 41555 35683
rect 41705 35649 41739 35683
rect 42809 35649 42843 35683
rect 43065 35649 43099 35683
rect 44833 35649 44867 35683
rect 46673 35649 46707 35683
rect 46949 35649 46983 35683
rect 24593 35581 24627 35615
rect 38761 35581 38795 35615
rect 39681 35581 39715 35615
rect 44649 35581 44683 35615
rect 27353 35445 27387 35479
rect 30573 35445 30607 35479
rect 34713 35445 34747 35479
rect 38301 35445 38335 35479
rect 40049 35445 40083 35479
rect 40509 35445 40543 35479
rect 44189 35445 44223 35479
rect 46673 35445 46707 35479
rect 26985 35241 27019 35275
rect 29009 35241 29043 35275
rect 32505 35241 32539 35275
rect 42901 35241 42935 35275
rect 44557 35241 44591 35275
rect 30113 35105 30147 35139
rect 30573 35105 30607 35139
rect 33517 35105 33551 35139
rect 44281 35105 44315 35139
rect 45477 35105 45511 35139
rect 45937 35105 45971 35139
rect 25605 35037 25639 35071
rect 25872 35037 25906 35071
rect 29193 35037 29227 35071
rect 29837 35037 29871 35071
rect 29929 35037 29963 35071
rect 30757 35037 30791 35071
rect 30941 35037 30975 35071
rect 31585 35037 31619 35071
rect 32689 35037 32723 35071
rect 33241 35037 33275 35071
rect 33333 35037 33367 35071
rect 37841 35037 37875 35071
rect 38577 35037 38611 35071
rect 40233 35037 40267 35071
rect 40417 35037 40451 35071
rect 40509 35037 40543 35071
rect 43177 35037 43211 35071
rect 43269 35037 43303 35071
rect 43361 35037 43395 35071
rect 43545 35037 43579 35071
rect 44189 35037 44223 35071
rect 45569 35037 45603 35071
rect 46949 35037 46983 35071
rect 47205 35037 47239 35071
rect 38853 34969 38887 35003
rect 31401 34901 31435 34935
rect 38025 34901 38059 34935
rect 40049 34901 40083 34935
rect 48329 34901 48363 34935
rect 25329 34697 25363 34731
rect 29653 34697 29687 34731
rect 35909 34697 35943 34731
rect 39681 34697 39715 34731
rect 43545 34697 43579 34731
rect 44465 34697 44499 34731
rect 47133 34697 47167 34731
rect 40877 34629 40911 34663
rect 44097 34629 44131 34663
rect 23949 34561 23983 34595
rect 24205 34561 24239 34595
rect 27261 34561 27295 34595
rect 27353 34561 27387 34595
rect 28273 34561 28307 34595
rect 28540 34561 28574 34595
rect 30389 34561 30423 34595
rect 30656 34561 30690 34595
rect 33701 34561 33735 34595
rect 33885 34561 33919 34595
rect 34529 34561 34563 34595
rect 34796 34561 34830 34595
rect 38209 34561 38243 34595
rect 38393 34561 38427 34595
rect 39497 34561 39531 34595
rect 39773 34561 39807 34595
rect 43177 34561 43211 34595
rect 43361 34561 43395 34595
rect 44281 34561 44315 34595
rect 44557 34561 44591 34595
rect 45845 34561 45879 34595
rect 46857 34561 46891 34595
rect 38577 34493 38611 34527
rect 39313 34493 39347 34527
rect 45937 34493 45971 34527
rect 47133 34493 47167 34527
rect 46213 34425 46247 34459
rect 27537 34357 27571 34391
rect 31769 34357 31803 34391
rect 34069 34357 34103 34391
rect 40969 34357 41003 34391
rect 46949 34357 46983 34391
rect 28917 34153 28951 34187
rect 35725 34153 35759 34187
rect 44005 34153 44039 34187
rect 48145 34153 48179 34187
rect 33701 34085 33735 34119
rect 38117 34085 38151 34119
rect 40049 34085 40083 34119
rect 30113 34017 30147 34051
rect 36737 34017 36771 34051
rect 40785 34017 40819 34051
rect 26065 33949 26099 33983
rect 29101 33949 29135 33983
rect 29837 33949 29871 33983
rect 29929 33949 29963 33983
rect 31217 33949 31251 33983
rect 34345 33949 34379 33983
rect 34897 33949 34931 33983
rect 35081 33949 35115 33983
rect 35265 33949 35299 33983
rect 35909 33949 35943 33983
rect 38761 33949 38795 33983
rect 38945 33949 38979 33983
rect 39037 33949 39071 33983
rect 40049 33949 40083 33983
rect 40233 33949 40267 33983
rect 40693 33949 40727 33983
rect 40877 33949 40911 33983
rect 44005 33949 44039 33983
rect 44189 33949 44223 33983
rect 48329 33949 48363 33983
rect 26332 33881 26366 33915
rect 30941 33881 30975 33915
rect 31309 33881 31343 33915
rect 33517 33881 33551 33915
rect 37004 33881 37038 33915
rect 27445 33813 27479 33847
rect 31125 33813 31159 33847
rect 31493 33813 31527 33847
rect 34161 33813 34195 33847
rect 38577 33813 38611 33847
rect 27169 33609 27203 33643
rect 35633 33609 35667 33643
rect 37473 33609 37507 33643
rect 38761 33609 38795 33643
rect 25237 33541 25271 33575
rect 30941 33541 30975 33575
rect 34520 33541 34554 33575
rect 36921 33541 36955 33575
rect 40969 33541 41003 33575
rect 24409 33473 24443 33507
rect 25053 33473 25087 33507
rect 27353 33473 27387 33507
rect 31217 33473 31251 33507
rect 33609 33473 33643 33507
rect 34253 33473 34287 33507
rect 36553 33473 36587 33507
rect 37749 33473 37783 33507
rect 37841 33473 37875 33507
rect 37933 33473 37967 33507
rect 38117 33473 38151 33507
rect 38577 33473 38611 33507
rect 38761 33473 38795 33507
rect 40785 33473 40819 33507
rect 41061 33473 41095 33507
rect 45293 33473 45327 33507
rect 24869 33405 24903 33439
rect 31125 33405 31159 33439
rect 33425 33405 33459 33439
rect 45201 33405 45235 33439
rect 2329 33269 2363 33303
rect 24225 33269 24259 33303
rect 31125 33269 31159 33303
rect 31401 33269 31435 33303
rect 33793 33269 33827 33303
rect 40785 33269 40819 33303
rect 45661 33269 45695 33303
rect 47961 33269 47995 33303
rect 45201 33065 45235 33099
rect 26709 32997 26743 33031
rect 1593 32929 1627 32963
rect 2789 32929 2823 32963
rect 32137 32929 32171 32963
rect 40509 32929 40543 32963
rect 40969 32929 41003 32963
rect 43453 32929 43487 32963
rect 43913 32929 43947 32963
rect 45385 32929 45419 32963
rect 45477 32929 45511 32963
rect 46489 32929 46523 32963
rect 24593 32861 24627 32895
rect 29929 32861 29963 32895
rect 31309 32861 31343 32895
rect 34161 32861 34195 32895
rect 36369 32861 36403 32895
rect 39129 32861 39163 32895
rect 39405 32861 39439 32895
rect 40601 32861 40635 32895
rect 41521 32861 41555 32895
rect 43545 32861 43579 32895
rect 44373 32871 44407 32905
rect 44557 32861 44591 32895
rect 45569 32861 45603 32895
rect 45661 32861 45695 32895
rect 1777 32793 1811 32827
rect 24860 32793 24894 32827
rect 26433 32793 26467 32827
rect 31493 32793 31527 32827
rect 32404 32793 32438 32827
rect 36636 32793 36670 32827
rect 41788 32793 41822 32827
rect 46673 32793 46707 32827
rect 48329 32793 48363 32827
rect 25973 32725 26007 32759
rect 26893 32725 26927 32759
rect 29745 32725 29779 32759
rect 31677 32725 31711 32759
rect 33517 32725 33551 32759
rect 33977 32725 34011 32759
rect 37749 32725 37783 32759
rect 38945 32725 38979 32759
rect 39313 32725 39347 32759
rect 42901 32725 42935 32759
rect 44557 32725 44591 32759
rect 2421 32521 2455 32555
rect 26341 32521 26375 32555
rect 30113 32521 30147 32555
rect 32321 32521 32355 32555
rect 41705 32521 41739 32555
rect 44833 32521 44867 32555
rect 47869 32521 47903 32555
rect 29000 32453 29034 32487
rect 32597 32453 32631 32487
rect 32807 32453 32841 32487
rect 42717 32453 42751 32487
rect 2329 32385 2363 32419
rect 25329 32385 25363 32419
rect 25973 32385 26007 32419
rect 28733 32385 28767 32419
rect 32505 32385 32539 32419
rect 32689 32385 32723 32419
rect 32965 32385 32999 32419
rect 37473 32385 37507 32419
rect 37657 32385 37691 32419
rect 37749 32385 37783 32419
rect 38945 32385 38979 32419
rect 40141 32385 40175 32419
rect 40969 32385 41003 32419
rect 41153 32385 41187 32419
rect 41521 32385 41555 32419
rect 42625 32385 42659 32419
rect 42809 32385 42843 32419
rect 43637 32385 43671 32419
rect 43821 32385 43855 32419
rect 43913 32385 43947 32419
rect 45293 32385 45327 32419
rect 46121 32385 46155 32419
rect 46949 32385 46983 32419
rect 47041 32385 47075 32419
rect 47777 32385 47811 32419
rect 25145 32317 25179 32351
rect 26249 32317 26283 32351
rect 26458 32317 26492 32351
rect 27169 32317 27203 32351
rect 39037 32317 39071 32351
rect 40234 32317 40268 32351
rect 40325 32317 40359 32351
rect 40417 32317 40451 32351
rect 41245 32317 41279 32351
rect 41337 32317 41371 32351
rect 45201 32317 45235 32351
rect 45477 32317 45511 32351
rect 46029 32317 46063 32351
rect 47225 32317 47259 32351
rect 27537 32249 27571 32283
rect 37473 32249 37507 32283
rect 39313 32249 39347 32283
rect 46489 32249 46523 32283
rect 25513 32181 25547 32215
rect 26617 32181 26651 32215
rect 27629 32181 27663 32215
rect 39957 32181 39991 32215
rect 43453 32181 43487 32215
rect 47133 32181 47167 32215
rect 30573 31977 30607 32011
rect 37381 31977 37415 32011
rect 38301 31977 38335 32011
rect 39405 31977 39439 32011
rect 40417 31977 40451 32011
rect 40877 31977 40911 32011
rect 44281 31977 44315 32011
rect 45201 31977 45235 32011
rect 48329 31977 48363 32011
rect 26157 31909 26191 31943
rect 45569 31909 45603 31943
rect 27169 31841 27203 31875
rect 34897 31841 34931 31875
rect 41061 31841 41095 31875
rect 41245 31841 41279 31875
rect 41337 31841 41371 31875
rect 45661 31841 45695 31875
rect 46949 31841 46983 31875
rect 26341 31773 26375 31807
rect 26617 31773 26651 31807
rect 27077 31773 27111 31807
rect 27261 31773 27295 31807
rect 27813 31773 27847 31807
rect 30205 31773 30239 31807
rect 30389 31773 30423 31807
rect 35081 31773 35115 31807
rect 35265 31773 35299 31807
rect 36093 31773 36127 31807
rect 38485 31773 38519 31807
rect 38669 31773 38703 31807
rect 38761 31773 38795 31807
rect 39313 31773 39347 31807
rect 39497 31773 39531 31807
rect 40049 31773 40083 31807
rect 41153 31773 41187 31807
rect 43913 31773 43947 31807
rect 45385 31773 45419 31807
rect 28058 31705 28092 31739
rect 40233 31705 40267 31739
rect 44097 31705 44131 31739
rect 47194 31705 47228 31739
rect 26525 31637 26559 31671
rect 29193 31637 29227 31671
rect 24869 31433 24903 31467
rect 28733 31433 28767 31467
rect 31769 31433 31803 31467
rect 32873 31433 32907 31467
rect 37565 31433 37599 31467
rect 40785 31433 40819 31467
rect 47041 31433 47075 31467
rect 29622 31365 29656 31399
rect 31309 31365 31343 31399
rect 32597 31365 32631 31399
rect 34314 31365 34348 31399
rect 46857 31365 46891 31399
rect 24133 31297 24167 31331
rect 24225 31297 24259 31331
rect 24409 31297 24443 31331
rect 25053 31297 25087 31331
rect 26249 31297 26283 31331
rect 26341 31297 26375 31331
rect 27169 31297 27203 31331
rect 27353 31297 27387 31331
rect 27445 31297 27479 31331
rect 27721 31297 27755 31331
rect 28917 31297 28951 31331
rect 31585 31297 31619 31331
rect 32321 31297 32355 31331
rect 32505 31297 32539 31331
rect 32689 31297 32723 31331
rect 36093 31297 36127 31331
rect 37473 31297 37507 31331
rect 38393 31297 38427 31331
rect 38485 31297 38519 31331
rect 38577 31297 38611 31331
rect 38761 31297 38795 31331
rect 40969 31297 41003 31331
rect 47133 31297 47167 31331
rect 26617 31229 26651 31263
rect 27537 31229 27571 31263
rect 29377 31229 29411 31263
rect 31493 31229 31527 31263
rect 34069 31229 34103 31263
rect 41153 31229 41187 31263
rect 41245 31229 41279 31263
rect 26525 31161 26559 31195
rect 46857 31161 46891 31195
rect 26065 31093 26099 31127
rect 27905 31093 27939 31127
rect 30757 31093 30791 31127
rect 31585 31093 31619 31127
rect 35449 31093 35483 31127
rect 35909 31093 35943 31127
rect 38117 31093 38151 31127
rect 30113 30889 30147 30923
rect 33609 30889 33643 30923
rect 38853 30889 38887 30923
rect 45845 30889 45879 30923
rect 29745 30753 29779 30787
rect 31217 30753 31251 30787
rect 40325 30753 40359 30787
rect 26525 30685 26559 30719
rect 26617 30685 26651 30719
rect 26801 30685 26835 30719
rect 26893 30685 26927 30719
rect 29929 30685 29963 30719
rect 31401 30685 31435 30719
rect 32229 30685 32263 30719
rect 34897 30685 34931 30719
rect 37473 30685 37507 30719
rect 37740 30685 37774 30719
rect 40509 30685 40543 30719
rect 40785 30685 40819 30719
rect 43177 30685 43211 30719
rect 43269 30685 43303 30719
rect 43361 30685 43395 30719
rect 43545 30685 43579 30719
rect 45201 30685 45235 30719
rect 45349 30685 45383 30719
rect 45666 30685 45700 30719
rect 46305 30685 46339 30719
rect 32496 30617 32530 30651
rect 35164 30617 35198 30651
rect 45477 30617 45511 30651
rect 45569 30617 45603 30651
rect 46397 30617 46431 30651
rect 26341 30549 26375 30583
rect 31585 30549 31619 30583
rect 36277 30549 36311 30583
rect 40693 30549 40727 30583
rect 42901 30549 42935 30583
rect 25421 30345 25455 30379
rect 33149 30345 33183 30379
rect 40141 30345 40175 30379
rect 41153 30345 41187 30379
rect 39129 30277 39163 30311
rect 39865 30277 39899 30311
rect 40877 30277 40911 30311
rect 43238 30277 43272 30311
rect 24297 30209 24331 30243
rect 31677 30209 31711 30243
rect 32321 30209 32355 30243
rect 32505 30209 32539 30243
rect 32689 30209 32723 30243
rect 33333 30209 33367 30243
rect 35357 30209 35391 30243
rect 35541 30209 35575 30243
rect 38853 30209 38887 30243
rect 39589 30209 39623 30243
rect 39773 30209 39807 30243
rect 39957 30209 39991 30243
rect 40601 30209 40635 30243
rect 40785 30209 40819 30243
rect 40969 30209 41003 30243
rect 44833 30209 44867 30243
rect 45017 30209 45051 30243
rect 45385 30209 45419 30243
rect 46029 30209 46063 30243
rect 47777 30209 47811 30243
rect 24041 30141 24075 30175
rect 39129 30141 39163 30175
rect 42993 30141 43027 30175
rect 45109 30141 45143 30175
rect 45201 30141 45235 30175
rect 46489 30141 46523 30175
rect 44373 30073 44407 30107
rect 31493 30005 31527 30039
rect 35357 30005 35391 30039
rect 38945 30005 38979 30039
rect 45569 30005 45603 30039
rect 46121 30005 46155 30039
rect 47225 30005 47259 30039
rect 47869 30005 47903 30039
rect 23397 29801 23431 29835
rect 28641 29801 28675 29835
rect 32689 29801 32723 29835
rect 39037 29801 39071 29835
rect 40049 29801 40083 29835
rect 40509 29801 40543 29835
rect 45753 29801 45787 29835
rect 22845 29733 22879 29767
rect 27261 29665 27295 29699
rect 35173 29665 35207 29699
rect 35265 29665 35299 29699
rect 42993 29665 43027 29699
rect 46489 29665 46523 29699
rect 22661 29597 22695 29631
rect 23673 29597 23707 29631
rect 23762 29597 23796 29631
rect 23857 29597 23891 29631
rect 24041 29597 24075 29631
rect 26341 29597 26375 29631
rect 26617 29597 26651 29631
rect 31309 29597 31343 29631
rect 31576 29597 31610 29631
rect 34897 29597 34931 29631
rect 36001 29597 36035 29631
rect 36185 29597 36219 29631
rect 38945 29597 38979 29631
rect 39129 29597 39163 29631
rect 40233 29597 40267 29631
rect 40325 29597 40359 29631
rect 40601 29597 40635 29631
rect 42717 29597 42751 29631
rect 42809 29597 42843 29631
rect 43085 29597 43119 29631
rect 43545 29597 43579 29631
rect 43729 29597 43763 29631
rect 43913 29597 43947 29631
rect 45661 29597 45695 29631
rect 27506 29529 27540 29563
rect 35382 29529 35416 29563
rect 43821 29529 43855 29563
rect 46673 29529 46707 29563
rect 48329 29529 48363 29563
rect 26157 29461 26191 29495
rect 26525 29461 26559 29495
rect 35541 29461 35575 29495
rect 36369 29461 36403 29495
rect 42533 29461 42567 29495
rect 44097 29461 44131 29495
rect 23305 29257 23339 29291
rect 23949 29257 23983 29291
rect 27169 29257 27203 29291
rect 40141 29257 40175 29291
rect 40785 29257 40819 29291
rect 41981 29257 42015 29291
rect 42901 29257 42935 29291
rect 43269 29257 43303 29291
rect 43913 29257 43947 29291
rect 34253 29189 34287 29223
rect 36185 29189 36219 29223
rect 24409 29121 24443 29155
rect 24593 29121 24627 29155
rect 26433 29121 26467 29155
rect 26617 29121 26651 29155
rect 27445 29121 27479 29155
rect 27537 29121 27571 29155
rect 27629 29121 27663 29155
rect 27813 29121 27847 29155
rect 28733 29121 28767 29155
rect 29000 29121 29034 29155
rect 30573 29121 30607 29155
rect 30757 29121 30791 29155
rect 35357 29121 35391 29155
rect 35449 29121 35483 29155
rect 35633 29121 35667 29155
rect 35725 29121 35759 29155
rect 37740 29121 37774 29155
rect 40049 29121 40083 29155
rect 40693 29121 40727 29155
rect 41889 29121 41923 29155
rect 43085 29121 43119 29155
rect 43361 29121 43395 29155
rect 43821 29121 43855 29155
rect 45825 29121 45859 29155
rect 23673 29053 23707 29087
rect 23765 29053 23799 29087
rect 31033 29053 31067 29087
rect 37473 29053 37507 29087
rect 45569 29053 45603 29087
rect 30941 28985 30975 29019
rect 34621 28985 34655 29019
rect 36461 28985 36495 29019
rect 38853 28985 38887 29019
rect 46949 28985 46983 29019
rect 24501 28917 24535 28951
rect 26433 28917 26467 28951
rect 30113 28917 30147 28951
rect 34713 28917 34747 28951
rect 35173 28917 35207 28951
rect 36645 28917 36679 28951
rect 47961 28917 47995 28951
rect 24961 28713 24995 28747
rect 26065 28713 26099 28747
rect 27813 28713 27847 28747
rect 29745 28713 29779 28747
rect 44097 28713 44131 28747
rect 45569 28713 45603 28747
rect 27261 28645 27295 28679
rect 40049 28645 40083 28679
rect 26801 28577 26835 28611
rect 35449 28577 35483 28611
rect 35541 28577 35575 28611
rect 41797 28577 41831 28611
rect 46029 28577 46063 28611
rect 46489 28577 46523 28611
rect 48237 28577 48271 28611
rect 23213 28509 23247 28543
rect 23489 28509 23523 28543
rect 24777 28509 24811 28543
rect 26065 28509 26099 28543
rect 26249 28509 26283 28543
rect 26893 28509 26927 28543
rect 27721 28509 27755 28543
rect 27905 28509 27939 28543
rect 30021 28509 30055 28543
rect 31217 28509 31251 28543
rect 35173 28509 35207 28543
rect 35357 28509 35391 28543
rect 35725 28509 35759 28543
rect 36553 28509 36587 28543
rect 36737 28509 36771 28543
rect 36829 28509 36863 28543
rect 40049 28509 40083 28543
rect 40233 28509 40267 28543
rect 40325 28509 40359 28543
rect 41521 28509 41555 28543
rect 41613 28509 41647 28543
rect 42257 28509 42291 28543
rect 42441 28509 42475 28543
rect 44005 28509 44039 28543
rect 45753 28509 45787 28543
rect 45937 28509 45971 28543
rect 24593 28441 24627 28475
rect 29745 28441 29779 28475
rect 31484 28441 31518 28475
rect 41797 28441 41831 28475
rect 46673 28441 46707 28475
rect 23029 28373 23063 28407
rect 23397 28373 23431 28407
rect 29929 28373 29963 28407
rect 32597 28373 32631 28407
rect 35909 28373 35943 28407
rect 36369 28373 36403 28407
rect 42349 28373 42383 28407
rect 33149 28169 33183 28203
rect 38025 28169 38059 28203
rect 39957 28169 39991 28203
rect 42073 28169 42107 28203
rect 45759 28169 45793 28203
rect 47869 28169 47903 28203
rect 24869 28101 24903 28135
rect 25085 28101 25119 28135
rect 26249 28101 26283 28135
rect 26617 28101 26651 28135
rect 32597 28101 32631 28135
rect 40960 28101 40994 28135
rect 45845 28101 45879 28135
rect 22937 28033 22971 28067
rect 23213 28033 23247 28067
rect 23673 28033 23707 28067
rect 23857 28033 23891 28067
rect 24041 28033 24075 28067
rect 24236 28033 24270 28067
rect 28641 28033 28675 28067
rect 30941 28033 30975 28067
rect 32321 28033 32355 28067
rect 33057 28033 33091 28067
rect 33241 28033 33275 28067
rect 35265 28033 35299 28067
rect 35357 28033 35391 28067
rect 35633 28033 35667 28067
rect 37933 28033 37967 28067
rect 38117 28033 38151 28067
rect 38844 28033 38878 28067
rect 40693 28033 40727 28067
rect 43168 28033 43202 28067
rect 45661 28033 45695 28067
rect 45937 28033 45971 28067
rect 46397 28033 46431 28067
rect 46581 28033 46615 28067
rect 47777 28033 47811 28067
rect 23958 27965 23992 27999
rect 31217 27965 31251 27999
rect 32597 27965 32631 27999
rect 35541 27965 35575 27999
rect 38577 27965 38611 27999
rect 42901 27965 42935 27999
rect 22753 27897 22787 27931
rect 25237 27897 25271 27931
rect 31033 27897 31067 27931
rect 23121 27829 23155 27863
rect 24409 27829 24443 27863
rect 25053 27829 25087 27863
rect 28733 27829 28767 27863
rect 31125 27829 31159 27863
rect 32413 27829 32447 27863
rect 35081 27829 35115 27863
rect 44281 27829 44315 27863
rect 46397 27829 46431 27863
rect 39129 27625 39163 27659
rect 40233 27625 40267 27659
rect 40417 27625 40451 27659
rect 42073 27625 42107 27659
rect 43177 27625 43211 27659
rect 43913 27625 43947 27659
rect 46121 27625 46155 27659
rect 46765 27625 46799 27659
rect 22753 27557 22787 27591
rect 26985 27557 27019 27591
rect 32137 27557 32171 27591
rect 39221 27557 39255 27591
rect 23581 27489 23615 27523
rect 23765 27489 23799 27523
rect 26525 27489 26559 27523
rect 29929 27489 29963 27523
rect 31769 27489 31803 27523
rect 39405 27489 39439 27523
rect 41705 27489 41739 27523
rect 45753 27489 45787 27523
rect 46673 27489 46707 27523
rect 46857 27489 46891 27523
rect 22661 27421 22695 27455
rect 22845 27421 22879 27455
rect 23489 27421 23523 27455
rect 23673 27421 23707 27455
rect 24593 27421 24627 27455
rect 24860 27421 24894 27455
rect 26617 27421 26651 27455
rect 27445 27421 27479 27455
rect 28089 27421 28123 27455
rect 31953 27421 31987 27455
rect 35081 27421 35115 27455
rect 35357 27421 35391 27455
rect 39129 27421 39163 27455
rect 41889 27421 41923 27455
rect 42993 27421 43027 27455
rect 43085 27421 43119 27455
rect 45937 27421 45971 27455
rect 46581 27421 46615 27455
rect 30196 27353 30230 27387
rect 33701 27353 33735 27387
rect 34897 27353 34931 27387
rect 40049 27353 40083 27387
rect 43269 27353 43303 27387
rect 43729 27353 43763 27387
rect 23305 27285 23339 27319
rect 25973 27285 26007 27319
rect 27537 27285 27571 27319
rect 28181 27285 28215 27319
rect 31309 27285 31343 27319
rect 33793 27285 33827 27319
rect 35265 27285 35299 27319
rect 40249 27285 40283 27319
rect 43929 27285 43963 27319
rect 44097 27285 44131 27319
rect 23397 27081 23431 27115
rect 25329 27081 25363 27115
rect 30113 27081 30147 27115
rect 31033 27081 31067 27115
rect 34345 27081 34379 27115
rect 34989 27081 35023 27115
rect 36921 27081 36955 27115
rect 43545 27081 43579 27115
rect 47225 27081 47259 27115
rect 30665 27013 30699 27047
rect 30881 27013 30915 27047
rect 43361 27013 43395 27047
rect 46112 27013 46146 27047
rect 23305 26945 23339 26979
rect 23489 26945 23523 26979
rect 25237 26945 25271 26979
rect 26065 26945 26099 26979
rect 27445 26945 27479 26979
rect 27538 26945 27572 26979
rect 27813 26945 27847 26979
rect 30021 26945 30055 26979
rect 30205 26945 30239 26979
rect 33232 26945 33266 26979
rect 34805 26945 34839 26979
rect 35081 26945 35115 26979
rect 35541 26945 35575 26979
rect 35808 26945 35842 26979
rect 43637 26945 43671 26979
rect 45845 26945 45879 26979
rect 47777 26945 47811 26979
rect 26157 26877 26191 26911
rect 32965 26877 32999 26911
rect 43361 26809 43395 26843
rect 26341 26741 26375 26775
rect 27261 26741 27295 26775
rect 27721 26741 27755 26775
rect 30849 26741 30883 26775
rect 34805 26741 34839 26775
rect 47869 26741 47903 26775
rect 32505 26537 32539 26571
rect 33517 26537 33551 26571
rect 33885 26537 33919 26571
rect 40417 26537 40451 26571
rect 43821 26537 43855 26571
rect 35725 26469 35759 26503
rect 39221 26469 39255 26503
rect 44373 26469 44407 26503
rect 35449 26401 35483 26435
rect 40509 26401 40543 26435
rect 46673 26401 46707 26435
rect 48237 26401 48271 26435
rect 26341 26333 26375 26367
rect 26525 26333 26559 26367
rect 26709 26333 26743 26367
rect 27169 26333 27203 26367
rect 27317 26333 27351 26367
rect 27445 26333 27479 26367
rect 27675 26333 27709 26367
rect 33701 26333 33735 26367
rect 33977 26333 34011 26367
rect 35357 26333 35391 26367
rect 38025 26333 38059 26367
rect 39497 26333 39531 26367
rect 40233 26333 40267 26367
rect 43637 26333 43671 26367
rect 43913 26333 43947 26367
rect 44557 26333 44591 26367
rect 44649 26333 44683 26367
rect 46489 26333 46523 26367
rect 27537 26265 27571 26299
rect 31217 26265 31251 26299
rect 36461 26265 36495 26299
rect 39221 26265 39255 26299
rect 39405 26265 39439 26299
rect 44373 26265 44407 26299
rect 27813 26197 27847 26231
rect 40049 26197 40083 26231
rect 43453 26197 43487 26231
rect 29929 25993 29963 26027
rect 35633 25993 35667 26027
rect 36185 25993 36219 26027
rect 40509 25993 40543 26027
rect 44649 25993 44683 26027
rect 28641 25925 28675 25959
rect 32413 25925 32447 25959
rect 37565 25925 37599 25959
rect 47225 25925 47259 25959
rect 22293 25857 22327 25891
rect 24297 25857 24331 25891
rect 27169 25857 27203 25891
rect 27353 25857 27387 25891
rect 27721 25857 27755 25891
rect 30849 25857 30883 25891
rect 31033 25857 31067 25891
rect 35541 25857 35575 25891
rect 35725 25857 35759 25891
rect 36461 25857 36495 25891
rect 36553 25857 36587 25891
rect 36645 25857 36679 25891
rect 36829 25857 36863 25891
rect 37473 25857 37507 25891
rect 37657 25857 37691 25891
rect 38301 25857 38335 25891
rect 39129 25857 39163 25891
rect 39396 25857 39430 25891
rect 43269 25857 43303 25891
rect 43536 25857 43570 25891
rect 47961 25857 47995 25891
rect 22201 25789 22235 25823
rect 24041 25789 24075 25823
rect 27445 25789 27479 25823
rect 27537 25789 27571 25823
rect 45385 25789 45419 25823
rect 45569 25789 45603 25823
rect 2329 25653 2363 25687
rect 22569 25653 22603 25687
rect 25421 25653 25455 25687
rect 27905 25653 27939 25687
rect 30849 25653 30883 25687
rect 32505 25653 32539 25687
rect 38393 25653 38427 25687
rect 23397 25449 23431 25483
rect 24685 25449 24719 25483
rect 28089 25449 28123 25483
rect 36369 25449 36403 25483
rect 38761 25381 38795 25415
rect 41429 25381 41463 25415
rect 1593 25313 1627 25347
rect 2789 25313 2823 25347
rect 31677 25313 31711 25347
rect 31861 25313 31895 25347
rect 46397 25313 46431 25347
rect 22753 25245 22787 25279
rect 23673 25245 23707 25279
rect 23765 25245 23799 25279
rect 23857 25245 23891 25279
rect 24041 25245 24075 25279
rect 24593 25245 24627 25279
rect 27445 25245 27479 25279
rect 27583 25245 27617 25279
rect 27910 25245 27944 25279
rect 29745 25245 29779 25279
rect 31585 25245 31619 25279
rect 35909 25245 35943 25279
rect 36369 25245 36403 25279
rect 36553 25245 36587 25279
rect 37013 25245 37047 25279
rect 37657 25245 37691 25279
rect 39037 25245 39071 25279
rect 41705 25245 41739 25279
rect 42165 25245 42199 25279
rect 42349 25245 42383 25279
rect 45937 25245 45971 25279
rect 1777 25177 1811 25211
rect 22569 25177 22603 25211
rect 27721 25177 27755 25211
rect 27813 25177 27847 25211
rect 29990 25177 30024 25211
rect 35541 25177 35575 25211
rect 38761 25177 38795 25211
rect 41429 25177 41463 25211
rect 46121 25177 46155 25211
rect 22937 25109 22971 25143
rect 31125 25109 31159 25143
rect 31861 25109 31895 25143
rect 37105 25109 37139 25143
rect 37749 25109 37783 25143
rect 38945 25109 38979 25143
rect 41613 25109 41647 25143
rect 42257 25109 42291 25143
rect 2421 24905 2455 24939
rect 23673 24905 23707 24939
rect 29837 24905 29871 24939
rect 31125 24905 31159 24939
rect 39865 24905 39899 24939
rect 41153 24905 41187 24939
rect 2329 24769 2363 24803
rect 22385 24769 22419 24803
rect 22569 24769 22603 24803
rect 23397 24769 23431 24803
rect 27629 24769 27663 24803
rect 27813 24769 27847 24803
rect 27905 24769 27939 24803
rect 28181 24769 28215 24803
rect 30021 24769 30055 24803
rect 30941 24769 30975 24803
rect 33425 24769 33459 24803
rect 33692 24769 33726 24803
rect 35265 24769 35299 24803
rect 35449 24769 35483 24803
rect 38752 24769 38786 24803
rect 40877 24769 40911 24803
rect 41797 24769 41831 24803
rect 42625 24769 42659 24803
rect 42892 24769 42926 24803
rect 46029 24769 46063 24803
rect 47041 24769 47075 24803
rect 47133 24769 47167 24803
rect 23029 24701 23063 24735
rect 23489 24701 23523 24735
rect 30297 24701 30331 24735
rect 30757 24701 30791 24735
rect 35725 24701 35759 24735
rect 38485 24701 38519 24735
rect 41153 24701 41187 24735
rect 41613 24701 41647 24735
rect 47961 24701 47995 24735
rect 22477 24633 22511 24667
rect 28089 24633 28123 24667
rect 30205 24633 30239 24667
rect 34805 24565 34839 24599
rect 35633 24565 35667 24599
rect 40969 24565 41003 24599
rect 41981 24565 42015 24599
rect 44005 24565 44039 24599
rect 46121 24565 46155 24599
rect 24961 24361 24995 24395
rect 28825 24361 28859 24395
rect 30021 24361 30055 24395
rect 32045 24361 32079 24395
rect 34897 24361 34931 24395
rect 36737 24361 36771 24395
rect 38669 24361 38703 24395
rect 42441 24361 42475 24395
rect 44649 24361 44683 24395
rect 45937 24361 45971 24395
rect 23305 24225 23339 24259
rect 23673 24225 23707 24259
rect 25053 24225 25087 24259
rect 32965 24225 32999 24259
rect 39037 24225 39071 24259
rect 42533 24225 42567 24259
rect 43269 24225 43303 24259
rect 2329 24157 2363 24191
rect 23765 24157 23799 24191
rect 24777 24157 24811 24191
rect 25513 24157 25547 24191
rect 25697 24157 25731 24191
rect 27169 24157 27203 24191
rect 27262 24157 27296 24191
rect 27445 24157 27479 24191
rect 27634 24157 27668 24191
rect 28549 24157 28583 24191
rect 28641 24157 28675 24191
rect 30665 24157 30699 24191
rect 34897 24157 34931 24191
rect 35173 24157 35207 24191
rect 36461 24157 36495 24191
rect 36553 24157 36587 24191
rect 36829 24157 36863 24191
rect 37473 24157 37507 24191
rect 37565 24157 37599 24191
rect 37749 24157 37783 24191
rect 37841 24157 37875 24191
rect 38853 24157 38887 24191
rect 39129 24157 39163 24191
rect 42257 24157 42291 24191
rect 45845 24157 45879 24191
rect 27537 24089 27571 24123
rect 29837 24089 29871 24123
rect 30053 24089 30087 24123
rect 30910 24089 30944 24123
rect 33232 24089 33266 24123
rect 42073 24089 42107 24123
rect 43514 24089 43548 24123
rect 23949 24021 23983 24055
rect 24593 24021 24627 24055
rect 25605 24021 25639 24055
rect 27813 24021 27847 24055
rect 30205 24021 30239 24055
rect 34345 24021 34379 24055
rect 35081 24021 35115 24055
rect 36277 24021 36311 24055
rect 37289 24021 37323 24055
rect 26249 23817 26283 23851
rect 30389 23817 30423 23851
rect 31141 23817 31175 23851
rect 31309 23817 31343 23851
rect 33793 23817 33827 23851
rect 38945 23817 38979 23851
rect 40157 23817 40191 23851
rect 40325 23817 40359 23851
rect 30941 23749 30975 23783
rect 36185 23749 36219 23783
rect 39957 23749 39991 23783
rect 41797 23749 41831 23783
rect 47225 23749 47259 23783
rect 2053 23681 2087 23715
rect 22293 23681 22327 23715
rect 23397 23681 23431 23715
rect 23489 23681 23523 23715
rect 23581 23681 23615 23715
rect 25237 23681 25271 23715
rect 25329 23681 25363 23715
rect 25513 23681 25547 23715
rect 26157 23681 26191 23715
rect 30297 23681 30331 23715
rect 30481 23681 30515 23715
rect 33701 23681 33735 23715
rect 33885 23681 33919 23715
rect 36001 23681 36035 23715
rect 36277 23681 36311 23715
rect 36369 23681 36403 23715
rect 37473 23681 37507 23715
rect 38853 23681 38887 23715
rect 41429 23681 41463 23715
rect 41522 23681 41556 23715
rect 41705 23681 41739 23715
rect 41935 23681 41969 23715
rect 2237 23613 2271 23647
rect 2789 23613 2823 23647
rect 22201 23613 22235 23647
rect 23305 23613 23339 23647
rect 25605 23613 25639 23647
rect 27721 23613 27755 23647
rect 27905 23613 27939 23647
rect 28549 23613 28583 23647
rect 37749 23613 37783 23647
rect 45385 23613 45419 23647
rect 45569 23613 45603 23647
rect 22661 23545 22695 23579
rect 23121 23477 23155 23511
rect 25605 23477 25639 23511
rect 31125 23477 31159 23511
rect 36553 23477 36587 23511
rect 37565 23477 37599 23511
rect 37657 23477 37691 23511
rect 40141 23477 40175 23511
rect 42073 23477 42107 23511
rect 2513 23273 2547 23307
rect 23489 23273 23523 23307
rect 26065 23273 26099 23307
rect 27997 23273 28031 23307
rect 28549 23273 28583 23307
rect 35081 23273 35115 23307
rect 45753 23273 45787 23307
rect 35265 23205 35299 23239
rect 40049 23205 40083 23239
rect 40877 23205 40911 23239
rect 23305 23137 23339 23171
rect 27537 23137 27571 23171
rect 28641 23137 28675 23171
rect 30849 23137 30883 23171
rect 36461 23137 36495 23171
rect 43269 23137 43303 23171
rect 44097 23137 44131 23171
rect 44189 23137 44223 23171
rect 2421 23069 2455 23103
rect 23213 23069 23247 23103
rect 24685 23069 24719 23103
rect 24952 23069 24986 23103
rect 26985 23069 27019 23103
rect 27077 23069 27111 23103
rect 27261 23069 27295 23103
rect 27445 23069 27479 23103
rect 28178 23069 28212 23103
rect 30573 23069 30607 23103
rect 30665 23069 30699 23103
rect 31309 23069 31343 23103
rect 36645 23069 36679 23103
rect 36921 23069 36955 23103
rect 37565 23069 37599 23103
rect 37841 23069 37875 23103
rect 38301 23069 38335 23103
rect 38485 23069 38519 23103
rect 40325 23069 40359 23103
rect 40785 23069 40819 23103
rect 41061 23069 41095 23103
rect 41613 23069 41647 23103
rect 43821 23069 43855 23103
rect 44005 23069 44039 23103
rect 44373 23069 44407 23103
rect 45661 23069 45695 23103
rect 46489 23069 46523 23103
rect 27353 23001 27387 23035
rect 31554 23001 31588 23035
rect 34897 23001 34931 23035
rect 35113 23001 35147 23035
rect 36829 23001 36863 23035
rect 40049 23001 40083 23035
rect 40233 23001 40267 23035
rect 46673 23001 46707 23035
rect 48329 23001 48363 23035
rect 28181 22933 28215 22967
rect 30573 22933 30607 22967
rect 32689 22933 32723 22967
rect 37381 22933 37415 22967
rect 37749 22933 37783 22967
rect 38393 22933 38427 22967
rect 40785 22933 40819 22967
rect 44557 22933 44591 22967
rect 27353 22729 27387 22763
rect 28457 22729 28491 22763
rect 36185 22729 36219 22763
rect 38117 22729 38151 22763
rect 39681 22729 39715 22763
rect 41521 22729 41555 22763
rect 43453 22729 43487 22763
rect 44281 22729 44315 22763
rect 47133 22729 47167 22763
rect 44189 22661 44223 22695
rect 44649 22661 44683 22695
rect 23213 22593 23247 22627
rect 23397 22593 23431 22627
rect 26433 22593 26467 22627
rect 27537 22593 27571 22627
rect 27629 22593 27663 22627
rect 27905 22593 27939 22627
rect 28365 22593 28399 22627
rect 29653 22593 29687 22627
rect 29837 22593 29871 22627
rect 30389 22593 30423 22627
rect 30573 22593 30607 22627
rect 30665 22593 30699 22627
rect 31217 22593 31251 22627
rect 31401 22593 31435 22627
rect 31493 22593 31527 22627
rect 33609 22593 33643 22627
rect 33876 22593 33910 22627
rect 36369 22593 36403 22627
rect 36461 22593 36495 22627
rect 36737 22593 36771 22627
rect 37565 22593 37599 22627
rect 37749 22593 37783 22627
rect 37841 22593 37875 22627
rect 37933 22593 37967 22627
rect 38945 22593 38979 22627
rect 39129 22593 39163 22627
rect 39313 22593 39347 22627
rect 39497 22593 39531 22627
rect 40141 22593 40175 22627
rect 40408 22593 40442 22627
rect 43361 22593 43395 22627
rect 44465 22593 44499 22627
rect 45109 22593 45143 22627
rect 47041 22593 47075 22627
rect 47961 22593 47995 22627
rect 29929 22525 29963 22559
rect 39221 22525 39255 22559
rect 44557 22525 44591 22559
rect 26525 22457 26559 22491
rect 27813 22457 27847 22491
rect 30389 22457 30423 22491
rect 31217 22457 31251 22491
rect 36645 22457 36679 22491
rect 45201 22457 45235 22491
rect 23213 22389 23247 22423
rect 29469 22389 29503 22423
rect 34989 22389 35023 22423
rect 31125 22185 31159 22219
rect 34069 22185 34103 22219
rect 42993 22185 43027 22219
rect 34161 22117 34195 22151
rect 34897 22117 34931 22151
rect 2789 22049 2823 22083
rect 23121 22049 23155 22083
rect 44005 22049 44039 22083
rect 1593 21981 1627 22015
rect 23305 21981 23339 22015
rect 23581 21981 23615 22015
rect 29745 21981 29779 22015
rect 34069 21981 34103 22015
rect 34897 21981 34931 22015
rect 35173 21981 35207 22015
rect 37289 21981 37323 22015
rect 40969 21981 41003 22015
rect 41153 21981 41187 22015
rect 41613 21981 41647 22015
rect 43913 21981 43947 22015
rect 46489 21981 46523 22015
rect 1777 21913 1811 21947
rect 29990 21913 30024 21947
rect 34345 21913 34379 21947
rect 35081 21913 35115 21947
rect 37556 21913 37590 21947
rect 41880 21913 41914 21947
rect 46673 21913 46707 21947
rect 48329 21913 48363 21947
rect 23489 21845 23523 21879
rect 38669 21845 38703 21879
rect 41061 21845 41095 21879
rect 44281 21845 44315 21879
rect 2881 21641 2915 21675
rect 22845 21641 22879 21675
rect 25789 21641 25823 21675
rect 30021 21641 30055 21675
rect 37841 21641 37875 21675
rect 44465 21641 44499 21675
rect 47133 21641 47167 21675
rect 29837 21573 29871 21607
rect 41613 21573 41647 21607
rect 42073 21573 42107 21607
rect 2329 21505 2363 21539
rect 2789 21505 2823 21539
rect 22569 21505 22603 21539
rect 22661 21505 22695 21539
rect 23535 21505 23569 21539
rect 23670 21508 23704 21542
rect 23765 21505 23799 21539
rect 23949 21505 23983 21539
rect 24409 21505 24443 21539
rect 24665 21505 24699 21539
rect 27537 21505 27571 21539
rect 27721 21505 27755 21539
rect 30113 21505 30147 21539
rect 37657 21505 37691 21539
rect 41705 21505 41739 21539
rect 41889 21505 41923 21539
rect 44097 21505 44131 21539
rect 47041 21505 47075 21539
rect 47961 21505 47995 21539
rect 37473 21437 37507 21471
rect 41981 21437 42015 21471
rect 44189 21437 44223 21471
rect 23305 21369 23339 21403
rect 27537 21301 27571 21335
rect 29837 21301 29871 21335
rect 24685 21097 24719 21131
rect 28273 21097 28307 21131
rect 31125 21097 31159 21131
rect 32965 21097 32999 21131
rect 44649 21097 44683 21131
rect 23213 20961 23247 20995
rect 25973 20961 26007 20995
rect 26893 20961 26927 20995
rect 43269 20961 43303 20995
rect 2329 20893 2363 20927
rect 23121 20893 23155 20927
rect 24593 20893 24627 20927
rect 24777 20893 24811 20927
rect 26065 20893 26099 20927
rect 29745 20893 29779 20927
rect 31585 20893 31619 20927
rect 34897 20893 34931 20927
rect 27160 20825 27194 20859
rect 29990 20825 30024 20859
rect 31852 20825 31886 20859
rect 35164 20825 35198 20859
rect 43514 20825 43548 20859
rect 23489 20757 23523 20791
rect 26433 20757 26467 20791
rect 36277 20757 36311 20791
rect 23305 20553 23339 20587
rect 26617 20553 26651 20587
rect 27261 20553 27295 20587
rect 28181 20553 28215 20587
rect 29745 20553 29779 20587
rect 31677 20553 31711 20587
rect 35357 20553 35391 20587
rect 42993 20553 43027 20587
rect 27169 20485 27203 20519
rect 2053 20417 2087 20451
rect 23213 20417 23247 20451
rect 23397 20417 23431 20451
rect 26249 20417 26283 20451
rect 27445 20417 27479 20451
rect 28089 20417 28123 20451
rect 29929 20417 29963 20451
rect 30205 20417 30239 20451
rect 31585 20417 31619 20451
rect 31769 20417 31803 20451
rect 32321 20417 32355 20451
rect 32588 20417 32622 20451
rect 34621 20417 34655 20451
rect 34805 20417 34839 20451
rect 34989 20417 35023 20451
rect 35173 20417 35207 20451
rect 35817 20417 35851 20451
rect 36001 20417 36035 20451
rect 36461 20417 36495 20451
rect 37749 20417 37783 20451
rect 38016 20417 38050 20451
rect 40509 20417 40543 20451
rect 40776 20417 40810 20451
rect 43269 20417 43303 20451
rect 43361 20417 43395 20451
rect 43453 20417 43487 20451
rect 43637 20417 43671 20451
rect 44097 20417 44131 20451
rect 44281 20417 44315 20451
rect 47041 20417 47075 20451
rect 2237 20349 2271 20383
rect 2789 20349 2823 20383
rect 26341 20349 26375 20383
rect 27537 20349 27571 20383
rect 30113 20349 30147 20383
rect 34897 20349 34931 20383
rect 35909 20281 35943 20315
rect 27537 20213 27571 20247
rect 33701 20213 33735 20247
rect 36553 20213 36587 20247
rect 39129 20213 39163 20247
rect 41889 20213 41923 20247
rect 44097 20213 44131 20247
rect 47133 20213 47167 20247
rect 47961 20213 47995 20247
rect 2513 20009 2547 20043
rect 32873 20009 32907 20043
rect 34161 20009 34195 20043
rect 34345 20009 34379 20043
rect 34897 20009 34931 20043
rect 37841 20009 37875 20043
rect 39037 20009 39071 20043
rect 41337 20009 41371 20043
rect 41981 20009 42015 20043
rect 43269 20009 43303 20043
rect 36277 19873 36311 19907
rect 40417 19873 40451 19907
rect 40509 19873 40543 19907
rect 43821 19873 43855 19907
rect 46489 19873 46523 19907
rect 46673 19873 46707 19907
rect 48237 19873 48271 19907
rect 2421 19805 2455 19839
rect 33149 19805 33183 19839
rect 33241 19805 33275 19839
rect 33333 19805 33367 19839
rect 33517 19805 33551 19839
rect 35081 19805 35115 19839
rect 35357 19805 35391 19839
rect 36001 19805 36035 19839
rect 36185 19805 36219 19839
rect 36737 19805 36771 19839
rect 38117 19805 38151 19839
rect 38209 19805 38243 19839
rect 38301 19805 38335 19839
rect 38485 19805 38519 19839
rect 38945 19805 38979 19839
rect 40233 19805 40267 19839
rect 41245 19805 41279 19839
rect 41337 19805 41371 19839
rect 41889 19805 41923 19839
rect 43177 19805 43211 19839
rect 43361 19805 43395 19839
rect 44005 19805 44039 19839
rect 33977 19737 34011 19771
rect 40969 19737 41003 19771
rect 34187 19669 34221 19703
rect 35265 19669 35299 19703
rect 35817 19669 35851 19703
rect 36829 19669 36863 19703
rect 40049 19669 40083 19703
rect 41061 19669 41095 19703
rect 44189 19669 44223 19703
rect 34161 19465 34195 19499
rect 37933 19465 37967 19499
rect 38577 19465 38611 19499
rect 40141 19465 40175 19499
rect 41245 19465 41279 19499
rect 43729 19465 43763 19499
rect 44557 19465 44591 19499
rect 35909 19397 35943 19431
rect 36093 19397 36127 19431
rect 32873 19329 32907 19363
rect 33057 19329 33091 19363
rect 33885 19329 33919 19363
rect 35082 19329 35116 19363
rect 35357 19329 35391 19363
rect 38301 19329 38335 19363
rect 39037 19329 39071 19363
rect 39405 19329 39439 19363
rect 39497 19329 39531 19363
rect 40601 19329 40635 19363
rect 41153 19329 41187 19363
rect 41337 19329 41371 19363
rect 43361 19329 43395 19363
rect 44373 19329 44407 19363
rect 44649 19329 44683 19363
rect 47041 19329 47075 19363
rect 32965 19261 32999 19295
rect 33517 19261 33551 19295
rect 33977 19261 34011 19295
rect 35173 19261 35207 19295
rect 35265 19261 35299 19295
rect 38393 19261 38427 19295
rect 40325 19261 40359 19295
rect 40417 19261 40451 19295
rect 40509 19261 40543 19295
rect 43269 19261 43303 19295
rect 44189 19261 44223 19295
rect 36277 19193 36311 19227
rect 34897 19125 34931 19159
rect 39681 19125 39715 19159
rect 47133 19125 47167 19159
rect 47961 19125 47995 19159
rect 34253 18921 34287 18955
rect 35725 18921 35759 18955
rect 38945 18921 38979 18955
rect 43821 18921 43855 18955
rect 40601 18853 40635 18887
rect 35541 18785 35575 18819
rect 37657 18785 37691 18819
rect 40141 18785 40175 18819
rect 46489 18785 46523 18819
rect 46673 18785 46707 18819
rect 48237 18785 48271 18819
rect 2329 18717 2363 18751
rect 34161 18717 34195 18751
rect 34345 18717 34379 18751
rect 35449 18717 35483 18751
rect 37749 18717 37783 18751
rect 38577 18717 38611 18751
rect 38761 18717 38795 18751
rect 40233 18717 40267 18751
rect 43821 18717 43855 18751
rect 44005 18717 44039 18751
rect 38117 18581 38151 18615
rect 35449 18377 35483 18411
rect 38577 18377 38611 18411
rect 40417 18377 40451 18411
rect 2053 18241 2087 18275
rect 35081 18241 35115 18275
rect 38485 18241 38519 18275
rect 38669 18241 38703 18275
rect 40049 18241 40083 18275
rect 47777 18241 47811 18275
rect 2237 18173 2271 18207
rect 2789 18173 2823 18207
rect 35173 18173 35207 18207
rect 40141 18173 40175 18207
rect 47869 18037 47903 18071
rect 2697 17833 2731 17867
rect 46673 17697 46707 17731
rect 48237 17697 48271 17731
rect 2605 17629 2639 17663
rect 46489 17629 46523 17663
rect 2237 17221 2271 17255
rect 47961 17153 47995 17187
rect 2053 17085 2087 17119
rect 2789 17085 2823 17119
rect 47225 16949 47259 16983
rect 2329 16745 2363 16779
rect 46489 16609 46523 16643
rect 48237 16609 48271 16643
rect 2789 16541 2823 16575
rect 2881 16473 2915 16507
rect 46673 16473 46707 16507
rect 47869 16201 47903 16235
rect 47777 16065 47811 16099
rect 1961 15453 1995 15487
rect 2421 15453 2455 15487
rect 47685 15453 47719 15487
rect 2513 15317 2547 15351
rect 2237 15045 2271 15079
rect 2053 14977 2087 15011
rect 47777 14977 47811 15011
rect 2789 14909 2823 14943
rect 47869 14773 47903 14807
rect 2789 14433 2823 14467
rect 46489 14433 46523 14467
rect 46673 14433 46707 14467
rect 48237 14433 48271 14467
rect 1593 14365 1627 14399
rect 1777 14297 1811 14331
rect 2881 14025 2915 14059
rect 2329 13889 2363 13923
rect 2789 13889 2823 13923
rect 47041 13889 47075 13923
rect 47133 13685 47167 13719
rect 47961 13685 47995 13719
rect 46489 13345 46523 13379
rect 46673 13345 46707 13379
rect 48237 13345 48271 13379
rect 47041 12801 47075 12835
rect 47133 12597 47167 12631
rect 47961 12597 47995 12631
rect 46489 12257 46523 12291
rect 46673 12257 46707 12291
rect 48237 12257 48271 12291
rect 2329 12189 2363 12223
rect 2053 11713 2087 11747
rect 47041 11713 47075 11747
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 47133 11509 47167 11543
rect 47961 11509 47995 11543
rect 2329 11305 2363 11339
rect 46489 11169 46523 11203
rect 46673 11169 46707 11203
rect 46949 11169 46983 11203
rect 2237 11101 2271 11135
rect 2329 10013 2363 10047
rect 2789 10013 2823 10047
rect 2881 9877 2915 9911
rect 2329 9605 2363 9639
rect 2145 9537 2179 9571
rect 2973 9469 3007 9503
rect 2145 8925 2179 8959
rect 2605 8925 2639 8959
rect 2697 8789 2731 8823
rect 2329 8517 2363 8551
rect 2145 8449 2179 8483
rect 41245 8449 41279 8483
rect 2789 8381 2823 8415
rect 41429 8381 41463 8415
rect 4077 7973 4111 8007
rect 1777 7905 1811 7939
rect 2973 7905 3007 7939
rect 47501 7905 47535 7939
rect 1593 7837 1627 7871
rect 3985 7837 4019 7871
rect 47777 7837 47811 7871
rect 2237 7429 2271 7463
rect 4537 7361 4571 7395
rect 2053 7293 2087 7327
rect 2789 7293 2823 7327
rect 5089 7293 5123 7327
rect 47961 7157 47995 7191
rect 2329 6953 2363 6987
rect 2973 6817 3007 6851
rect 4077 6817 4111 6851
rect 46489 6817 46523 6851
rect 48237 6817 48271 6851
rect 3985 6749 4019 6783
rect 46673 6681 46707 6715
rect 47869 6409 47903 6443
rect 46397 6273 46431 6307
rect 47041 6273 47075 6307
rect 47777 6273 47811 6307
rect 2145 6205 2179 6239
rect 2329 6205 2363 6239
rect 2973 6205 3007 6239
rect 4629 6069 4663 6103
rect 46489 6069 46523 6103
rect 47133 6069 47167 6103
rect 2329 5865 2363 5899
rect 2881 5865 2915 5899
rect 5457 5729 5491 5763
rect 46673 5729 46707 5763
rect 48237 5729 48271 5763
rect 2789 5661 2823 5695
rect 3985 5661 4019 5695
rect 4813 5661 4847 5695
rect 46029 5661 46063 5695
rect 46489 5661 46523 5695
rect 4077 5525 4111 5559
rect 2329 5253 2363 5287
rect 2145 5185 2179 5219
rect 4445 5185 4479 5219
rect 5181 5185 5215 5219
rect 5825 5185 5859 5219
rect 45385 5185 45419 5219
rect 47961 5185 47995 5219
rect 2789 5117 2823 5151
rect 45569 5117 45603 5151
rect 47225 5117 47259 5151
rect 4537 4981 4571 5015
rect 5273 4981 5307 5015
rect 5917 4981 5951 5015
rect 44925 4981 44959 5015
rect 44557 4777 44591 4811
rect 2973 4641 3007 4675
rect 4905 4641 4939 4675
rect 5549 4641 5583 4675
rect 46489 4641 46523 4675
rect 1593 4573 1627 4607
rect 4261 4573 4295 4607
rect 4721 4573 4755 4607
rect 7205 4573 7239 4607
rect 40233 4573 40267 4607
rect 44465 4573 44499 4607
rect 45201 4573 45235 4607
rect 45845 4573 45879 4607
rect 1777 4505 1811 4539
rect 46673 4505 46707 4539
rect 48329 4505 48363 4539
rect 45293 4437 45327 4471
rect 45937 4437 45971 4471
rect 2605 4233 2639 4267
rect 2053 4097 2087 4131
rect 2513 4097 2547 4131
rect 3157 4097 3191 4131
rect 7021 4097 7055 4131
rect 8309 4097 8343 4131
rect 10425 4097 10459 4131
rect 13001 4097 13035 4131
rect 43729 4097 43763 4131
rect 44373 4097 44407 4131
rect 47961 4097 47995 4131
rect 3801 4029 3835 4063
rect 3985 4029 4019 4063
rect 4261 4029 4295 4063
rect 38669 4029 38703 4063
rect 38853 4029 38887 4063
rect 39497 4029 39531 4063
rect 45385 4029 45419 4063
rect 45569 4029 45603 4063
rect 47225 4029 47259 4063
rect 3249 3893 3283 3927
rect 7113 3893 7147 3927
rect 7849 3893 7883 3927
rect 8401 3893 8435 3927
rect 10517 3893 10551 3927
rect 12449 3893 12483 3927
rect 13093 3893 13127 3927
rect 25421 3893 25455 3927
rect 26157 3893 26191 3927
rect 41153 3893 41187 3927
rect 41797 3893 41831 3927
rect 43821 3893 43855 3927
rect 44465 3893 44499 3927
rect 1593 3553 1627 3587
rect 1777 3553 1811 3587
rect 2789 3553 2823 3587
rect 5089 3553 5123 3587
rect 6193 3553 6227 3587
rect 6653 3553 6687 3587
rect 10517 3553 10551 3587
rect 10977 3553 11011 3587
rect 25881 3553 25915 3587
rect 26433 3553 26467 3587
rect 39405 3553 39439 3587
rect 40509 3553 40543 3587
rect 41245 3553 41279 3587
rect 45661 3553 45695 3587
rect 48145 3553 48179 3587
rect 4445 3485 4479 3519
rect 5549 3485 5583 3519
rect 10333 3485 10367 3519
rect 13185 3485 13219 3519
rect 16957 3485 16991 3519
rect 17417 3485 17451 3519
rect 18889 3485 18923 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 20729 3485 20763 3519
rect 22201 3485 22235 3519
rect 22661 3485 22695 3519
rect 24593 3485 24627 3519
rect 25237 3485 25271 3519
rect 28365 3485 28399 3519
rect 31861 3485 31895 3519
rect 32321 3485 32355 3519
rect 38025 3485 38059 3519
rect 38853 3485 38887 3519
rect 39313 3485 39347 3519
rect 42809 3485 42843 3519
rect 43913 3485 43947 3519
rect 44557 3485 44591 3519
rect 5641 3417 5675 3451
rect 6377 3417 6411 3451
rect 25329 3417 25363 3451
rect 26065 3417 26099 3451
rect 40693 3417 40727 3451
rect 45845 3417 45879 3451
rect 47501 3417 47535 3451
rect 17509 3349 17543 3383
rect 19533 3349 19567 3383
rect 20821 3349 20855 3383
rect 22753 3349 22787 3383
rect 24685 3349 24719 3383
rect 32413 3349 32447 3383
rect 38117 3349 38151 3383
rect 42901 3349 42935 3383
rect 4353 3077 4387 3111
rect 7757 3077 7791 3111
rect 13185 3077 13219 3111
rect 17049 3077 17083 3111
rect 19809 3077 19843 3111
rect 22201 3077 22235 3111
rect 24961 3077 24995 3111
rect 32505 3077 32539 3111
rect 38577 3077 38611 3111
rect 41429 3077 41463 3111
rect 42809 3077 42843 3111
rect 45109 3077 45143 3111
rect 1869 3009 1903 3043
rect 4169 3009 4203 3043
rect 7573 3009 7607 3043
rect 10517 3009 10551 3043
rect 12357 3009 12391 3043
rect 13001 3009 13035 3043
rect 16865 3009 16899 3043
rect 22017 3009 22051 3043
rect 24777 3009 24811 3043
rect 27445 3009 27479 3043
rect 32321 3009 32355 3043
rect 38393 3009 38427 3043
rect 40693 3009 40727 3043
rect 41337 3009 41371 3043
rect 42625 3009 42659 3043
rect 44925 3009 44959 3043
rect 47961 3009 47995 3043
rect 2053 2941 2087 2975
rect 2881 2941 2915 2975
rect 5181 2941 5215 2975
rect 8033 2941 8067 2975
rect 13553 2941 13587 2975
rect 17417 2941 17451 2975
rect 19625 2941 19659 2975
rect 20637 2941 20671 2975
rect 22569 2941 22603 2975
rect 25789 2941 25823 2975
rect 27629 2941 27663 2975
rect 27905 2941 27939 2975
rect 32781 2941 32815 2975
rect 40233 2941 40267 2975
rect 43085 2941 43119 2975
rect 45385 2941 45419 2975
rect 7113 2805 7147 2839
rect 12449 2805 12483 2839
rect 40785 2805 40819 2839
rect 4169 2601 4203 2635
rect 4721 2601 4755 2635
rect 5641 2601 5675 2635
rect 27629 2601 27663 2635
rect 38945 2601 38979 2635
rect 47869 2601 47903 2635
rect 2053 2465 2087 2499
rect 6745 2465 6779 2499
rect 7205 2465 7239 2499
rect 11897 2465 11931 2499
rect 12081 2465 12115 2499
rect 12909 2465 12943 2499
rect 19625 2465 19659 2499
rect 19901 2465 19935 2499
rect 24869 2465 24903 2499
rect 40049 2465 40083 2499
rect 40233 2465 40267 2499
rect 40601 2465 40635 2499
rect 42809 2465 42843 2499
rect 42993 2465 43027 2499
rect 45201 2465 45235 2499
rect 45385 2465 45419 2499
rect 45753 2465 45787 2499
rect 1593 2397 1627 2431
rect 4629 2397 4663 2431
rect 5549 2397 5583 2431
rect 19441 2397 19475 2431
rect 24593 2397 24627 2431
rect 27537 2397 27571 2431
rect 47777 2397 47811 2431
rect 1777 2329 1811 2363
rect 6929 2329 6963 2363
rect 44649 2329 44683 2363
<< metal1 >>
rect 14 48764 20 48816
rect 72 48804 78 48816
rect 8018 48804 8024 48816
rect 72 48776 8024 48804
rect 72 48764 78 48776
rect 8018 48764 8024 48776
rect 8076 48764 8082 48816
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 4890 47172 4896 47184
rect 2056 47144 4896 47172
rect 2056 47048 2084 47144
rect 4890 47132 4896 47144
rect 4948 47132 4954 47184
rect 3510 47064 3516 47116
rect 3568 47104 3574 47116
rect 7006 47104 7012 47116
rect 3568 47076 7012 47104
rect 3568 47064 3574 47076
rect 7006 47064 7012 47076
rect 7064 47064 7070 47116
rect 47210 47104 47216 47116
rect 47171 47076 47216 47104
rect 47210 47064 47216 47076
rect 47268 47064 47274 47116
rect 1949 47039 2007 47045
rect 1949 47005 1961 47039
rect 1995 47036 2007 47039
rect 2038 47036 2044 47048
rect 1995 47008 2044 47036
rect 1995 47005 2007 47008
rect 1949 46999 2007 47005
rect 2038 46996 2044 47008
rect 2096 46996 2102 47048
rect 2682 47036 2688 47048
rect 2643 47008 2688 47036
rect 2682 46996 2688 47008
rect 2740 46996 2746 47048
rect 4154 46996 4160 47048
rect 4212 47036 4218 47048
rect 4525 47039 4583 47045
rect 4525 47036 4537 47039
rect 4212 47008 4537 47036
rect 4212 46996 4218 47008
rect 4525 47005 4537 47008
rect 4571 47005 4583 47039
rect 4525 46999 4583 47005
rect 5169 47039 5227 47045
rect 5169 47005 5181 47039
rect 5215 47036 5227 47039
rect 5534 47036 5540 47048
rect 5215 47008 5540 47036
rect 5215 47005 5227 47008
rect 5169 46999 5227 47005
rect 5534 46996 5540 47008
rect 5592 46996 5598 47048
rect 5629 47039 5687 47045
rect 5629 47005 5641 47039
rect 5675 47036 5687 47039
rect 5718 47036 5724 47048
rect 5675 47008 5724 47036
rect 5675 47005 5687 47008
rect 5629 46999 5687 47005
rect 5718 46996 5724 47008
rect 5776 46996 5782 47048
rect 6546 46996 6552 47048
rect 6604 47036 6610 47048
rect 6733 47039 6791 47045
rect 6733 47036 6745 47039
rect 6604 47008 6745 47036
rect 6604 46996 6610 47008
rect 6733 47005 6745 47008
rect 6779 47005 6791 47039
rect 7374 47036 7380 47048
rect 7335 47008 7380 47036
rect 6733 46999 6791 47005
rect 7374 46996 7380 47008
rect 7432 46996 7438 47048
rect 8018 47036 8024 47048
rect 7979 47008 8024 47036
rect 8018 46996 8024 47008
rect 8076 46996 8082 47048
rect 8386 46996 8392 47048
rect 8444 47036 8450 47048
rect 9309 47039 9367 47045
rect 9309 47036 9321 47039
rect 8444 47008 9321 47036
rect 8444 46996 8450 47008
rect 9309 47005 9321 47008
rect 9355 47005 9367 47039
rect 12526 47036 12532 47048
rect 12487 47008 12532 47036
rect 9309 46999 9367 47005
rect 12526 46996 12532 47008
rect 12584 46996 12590 47048
rect 14550 47036 14556 47048
rect 14511 47008 14556 47036
rect 14550 46996 14556 47008
rect 14608 46996 14614 47048
rect 15194 47036 15200 47048
rect 15155 47008 15200 47036
rect 15194 46996 15200 47008
rect 15252 46996 15258 47048
rect 22462 46996 22468 47048
rect 22520 47036 22526 47048
rect 23017 47039 23075 47045
rect 23017 47036 23029 47039
rect 22520 47008 23029 47036
rect 22520 46996 22526 47008
rect 23017 47005 23029 47008
rect 23063 47005 23075 47039
rect 25314 47036 25320 47048
rect 25275 47008 25320 47036
rect 23017 46999 23075 47005
rect 25314 46996 25320 47008
rect 25372 46996 25378 47048
rect 27154 46996 27160 47048
rect 27212 47036 27218 47048
rect 27341 47039 27399 47045
rect 27341 47036 27353 47039
rect 27212 47008 27353 47036
rect 27212 46996 27218 47008
rect 27341 47005 27353 47008
rect 27387 47005 27399 47039
rect 27982 47036 27988 47048
rect 27943 47008 27988 47036
rect 27341 46999 27399 47005
rect 27982 46996 27988 47008
rect 28040 46996 28046 47048
rect 29086 47036 29092 47048
rect 29047 47008 29092 47036
rect 29086 46996 29092 47008
rect 29144 46996 29150 47048
rect 29914 47036 29920 47048
rect 29875 47008 29920 47036
rect 29914 46996 29920 47008
rect 29972 46996 29978 47048
rect 33226 47036 33232 47048
rect 33187 47008 33232 47036
rect 33226 46996 33232 47008
rect 33284 46996 33290 47048
rect 38289 47039 38347 47045
rect 38289 47005 38301 47039
rect 38335 47036 38347 47039
rect 39758 47036 39764 47048
rect 38335 47008 39764 47036
rect 38335 47005 38347 47008
rect 38289 46999 38347 47005
rect 39758 46996 39764 47008
rect 39816 46996 39822 47048
rect 41601 47039 41659 47045
rect 41601 47005 41613 47039
rect 41647 47036 41659 47039
rect 42610 47036 42616 47048
rect 41647 47008 42616 47036
rect 41647 47005 41659 47008
rect 41601 46999 41659 47005
rect 42610 46996 42616 47008
rect 42668 46996 42674 47048
rect 44634 47036 44640 47048
rect 44595 47008 44640 47036
rect 44634 46996 44640 47008
rect 44692 46996 44698 47048
rect 45370 47036 45376 47048
rect 45331 47008 45376 47036
rect 45370 46996 45376 47008
rect 45428 46996 45434 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 3237 46971 3295 46977
rect 3237 46937 3249 46971
rect 3283 46968 3295 46971
rect 4798 46968 4804 46980
rect 3283 46940 4804 46968
rect 3283 46937 3295 46940
rect 3237 46931 3295 46937
rect 4798 46928 4804 46940
rect 4856 46928 4862 46980
rect 45554 46928 45560 46980
rect 45612 46968 45618 46980
rect 47854 46968 47860 46980
rect 45612 46940 45657 46968
rect 47815 46940 47860 46968
rect 45612 46928 45618 46940
rect 47854 46928 47860 46940
rect 47912 46928 47918 46980
rect 1762 46860 1768 46912
rect 1820 46900 1826 46912
rect 2041 46903 2099 46909
rect 2041 46900 2053 46903
rect 1820 46872 2053 46900
rect 1820 46860 1826 46872
rect 2041 46869 2053 46872
rect 2087 46869 2099 46903
rect 2041 46863 2099 46869
rect 5721 46903 5779 46909
rect 5721 46869 5733 46903
rect 5767 46900 5779 46903
rect 6730 46900 6736 46912
rect 5767 46872 6736 46900
rect 5767 46869 5779 46872
rect 5721 46863 5779 46869
rect 6730 46860 6736 46872
rect 6788 46860 6794 46912
rect 7834 46900 7840 46912
rect 7795 46872 7840 46900
rect 7834 46860 7840 46872
rect 7892 46860 7898 46912
rect 9122 46900 9128 46912
rect 9083 46872 9128 46900
rect 9122 46860 9128 46872
rect 9180 46860 9186 46912
rect 27798 46900 27804 46912
rect 27759 46872 27804 46900
rect 27798 46860 27804 46872
rect 27856 46860 27862 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 7374 46696 7380 46708
rect 1872 46668 7380 46696
rect 1872 46569 1900 46668
rect 7374 46656 7380 46668
rect 7432 46656 7438 46708
rect 2041 46631 2099 46637
rect 2041 46597 2053 46631
rect 2087 46628 2099 46631
rect 4062 46628 4068 46640
rect 2087 46600 4068 46628
rect 2087 46597 2099 46600
rect 2041 46591 2099 46597
rect 4062 46588 4068 46600
rect 4120 46588 4126 46640
rect 6730 46628 6736 46640
rect 6691 46600 6736 46628
rect 6730 46588 6736 46600
rect 6788 46588 6794 46640
rect 12526 46628 12532 46640
rect 12176 46600 12532 46628
rect 1857 46563 1915 46569
rect 1857 46529 1869 46563
rect 1903 46529 1915 46563
rect 4154 46560 4160 46572
rect 4115 46532 4160 46560
rect 1857 46523 1915 46529
rect 4154 46520 4160 46532
rect 4212 46520 4218 46572
rect 6546 46560 6552 46572
rect 6507 46532 6552 46560
rect 6546 46520 6552 46532
rect 6604 46520 6610 46572
rect 12176 46569 12204 46600
rect 12526 46588 12532 46600
rect 12584 46588 12590 46640
rect 15194 46628 15200 46640
rect 14476 46600 15200 46628
rect 14476 46569 14504 46600
rect 15194 46588 15200 46600
rect 15252 46588 15258 46640
rect 25314 46628 25320 46640
rect 24780 46600 25320 46628
rect 12161 46563 12219 46569
rect 12161 46529 12173 46563
rect 12207 46529 12219 46563
rect 12161 46523 12219 46529
rect 14461 46563 14519 46569
rect 14461 46529 14473 46563
rect 14507 46529 14519 46563
rect 22462 46560 22468 46572
rect 22423 46532 22468 46560
rect 14461 46523 14519 46529
rect 22462 46520 22468 46532
rect 22520 46520 22526 46572
rect 24780 46569 24808 46600
rect 25314 46588 25320 46600
rect 25372 46588 25378 46640
rect 33226 46628 33232 46640
rect 32968 46600 33232 46628
rect 24765 46563 24823 46569
rect 24765 46529 24777 46563
rect 24811 46529 24823 46563
rect 27154 46560 27160 46572
rect 27115 46532 27160 46560
rect 24765 46523 24823 46529
rect 27154 46520 27160 46532
rect 27212 46520 27218 46572
rect 29086 46520 29092 46572
rect 29144 46560 29150 46572
rect 32968 46569 32996 46600
rect 33226 46588 33232 46600
rect 33284 46588 33290 46640
rect 47213 46631 47271 46637
rect 47213 46597 47225 46631
rect 47259 46628 47271 46631
rect 48314 46628 48320 46640
rect 47259 46600 48320 46628
rect 47259 46597 47271 46600
rect 47213 46591 47271 46597
rect 48314 46588 48320 46600
rect 48372 46588 48378 46640
rect 29457 46563 29515 46569
rect 29457 46560 29469 46563
rect 29144 46532 29469 46560
rect 29144 46520 29150 46532
rect 29457 46529 29469 46532
rect 29503 46529 29515 46563
rect 29457 46523 29515 46529
rect 32953 46563 33011 46569
rect 32953 46529 32965 46563
rect 32999 46529 33011 46563
rect 39758 46560 39764 46572
rect 39719 46532 39764 46560
rect 32953 46523 33011 46529
rect 39758 46520 39764 46532
rect 39816 46520 39822 46572
rect 42610 46560 42616 46572
rect 42571 46532 42616 46560
rect 42610 46520 42616 46532
rect 42668 46520 42674 46572
rect 44634 46520 44640 46572
rect 44692 46560 44698 46572
rect 45373 46563 45431 46569
rect 45373 46560 45385 46563
rect 44692 46532 45385 46560
rect 44692 46520 44698 46532
rect 45373 46529 45385 46532
rect 45419 46529 45431 46563
rect 45373 46523 45431 46529
rect 2590 46452 2596 46504
rect 2648 46492 2654 46504
rect 2777 46495 2835 46501
rect 2777 46492 2789 46495
rect 2648 46464 2789 46492
rect 2648 46452 2654 46464
rect 2777 46461 2789 46464
rect 2823 46461 2835 46495
rect 2777 46455 2835 46461
rect 4341 46495 4399 46501
rect 4341 46461 4353 46495
rect 4387 46492 4399 46495
rect 4614 46492 4620 46504
rect 4387 46464 4620 46492
rect 4387 46461 4399 46464
rect 4341 46455 4399 46461
rect 4614 46452 4620 46464
rect 4672 46452 4678 46504
rect 4706 46452 4712 46504
rect 4764 46492 4770 46504
rect 7006 46492 7012 46504
rect 4764 46464 4809 46492
rect 6967 46464 7012 46492
rect 4764 46452 4770 46464
rect 7006 46452 7012 46464
rect 7064 46452 7070 46504
rect 12345 46495 12403 46501
rect 12345 46461 12357 46495
rect 12391 46492 12403 46495
rect 12434 46492 12440 46504
rect 12391 46464 12440 46492
rect 12391 46461 12403 46464
rect 12345 46455 12403 46461
rect 12434 46452 12440 46464
rect 12492 46452 12498 46504
rect 12894 46492 12900 46504
rect 12855 46464 12900 46492
rect 12894 46452 12900 46464
rect 12952 46452 12958 46504
rect 14642 46492 14648 46504
rect 14603 46464 14648 46492
rect 14642 46452 14648 46464
rect 14700 46452 14706 46504
rect 15470 46492 15476 46504
rect 15431 46464 15476 46492
rect 15470 46452 15476 46464
rect 15528 46452 15534 46504
rect 22649 46495 22707 46501
rect 22649 46461 22661 46495
rect 22695 46492 22707 46495
rect 22922 46492 22928 46504
rect 22695 46464 22928 46492
rect 22695 46461 22707 46464
rect 22649 46455 22707 46461
rect 22922 46452 22928 46464
rect 22980 46452 22986 46504
rect 23198 46492 23204 46504
rect 23159 46464 23204 46492
rect 23198 46452 23204 46464
rect 23256 46452 23262 46504
rect 24946 46492 24952 46504
rect 24907 46464 24952 46492
rect 24946 46452 24952 46464
rect 25004 46452 25010 46504
rect 25774 46492 25780 46504
rect 25735 46464 25780 46492
rect 25774 46452 25780 46464
rect 25832 46452 25838 46504
rect 26970 46452 26976 46504
rect 27028 46492 27034 46504
rect 27341 46495 27399 46501
rect 27341 46492 27353 46495
rect 27028 46464 27353 46492
rect 27028 46452 27034 46464
rect 27341 46461 27353 46464
rect 27387 46461 27399 46495
rect 27341 46455 27399 46461
rect 27617 46495 27675 46501
rect 27617 46461 27629 46495
rect 27663 46461 27675 46495
rect 29638 46492 29644 46504
rect 29599 46464 29644 46492
rect 27617 46455 27675 46461
rect 1946 46384 1952 46436
rect 2004 46424 2010 46436
rect 2958 46424 2964 46436
rect 2004 46396 2964 46424
rect 2004 46384 2010 46396
rect 2958 46384 2964 46396
rect 3016 46384 3022 46436
rect 27062 46384 27068 46436
rect 27120 46424 27126 46436
rect 27632 46424 27660 46455
rect 29638 46452 29644 46464
rect 29696 46452 29702 46504
rect 29730 46452 29736 46504
rect 29788 46492 29794 46504
rect 29917 46495 29975 46501
rect 29917 46492 29929 46495
rect 29788 46464 29929 46492
rect 29788 46452 29794 46464
rect 29917 46461 29929 46464
rect 29963 46461 29975 46495
rect 29917 46455 29975 46461
rect 33137 46495 33195 46501
rect 33137 46461 33149 46495
rect 33183 46492 33195 46495
rect 33226 46492 33232 46504
rect 33183 46464 33232 46492
rect 33183 46461 33195 46464
rect 33137 46455 33195 46461
rect 33226 46452 33232 46464
rect 33284 46452 33290 46504
rect 33502 46492 33508 46504
rect 33463 46464 33508 46492
rect 33502 46452 33508 46464
rect 33560 46452 33566 46504
rect 36541 46495 36599 46501
rect 36541 46461 36553 46495
rect 36587 46492 36599 46495
rect 37461 46495 37519 46501
rect 37461 46492 37473 46495
rect 36587 46464 37473 46492
rect 36587 46461 36599 46464
rect 36541 46455 36599 46461
rect 37461 46461 37473 46464
rect 37507 46461 37519 46495
rect 37642 46492 37648 46504
rect 37603 46464 37648 46492
rect 37461 46455 37519 46461
rect 37642 46452 37648 46464
rect 37700 46452 37706 46504
rect 37921 46495 37979 46501
rect 37921 46461 37933 46495
rect 37967 46461 37979 46495
rect 39942 46492 39948 46504
rect 39903 46464 39948 46492
rect 37921 46455 37979 46461
rect 27120 46396 27660 46424
rect 27120 46384 27126 46396
rect 36722 46384 36728 46436
rect 36780 46424 36786 46436
rect 37936 46424 37964 46455
rect 39942 46452 39948 46464
rect 40000 46452 40006 46504
rect 40221 46495 40279 46501
rect 40221 46461 40233 46495
rect 40267 46461 40279 46495
rect 42794 46492 42800 46504
rect 42755 46464 42800 46492
rect 40221 46455 40279 46461
rect 36780 46396 37964 46424
rect 36780 46384 36786 46396
rect 38654 46384 38660 46436
rect 38712 46424 38718 46436
rect 40236 46424 40264 46455
rect 42794 46452 42800 46464
rect 42852 46452 42858 46504
rect 43073 46495 43131 46501
rect 43073 46461 43085 46495
rect 43119 46461 43131 46495
rect 43073 46455 43131 46461
rect 45557 46495 45615 46501
rect 45557 46461 45569 46495
rect 45603 46492 45615 46495
rect 48038 46492 48044 46504
rect 45603 46464 48044 46492
rect 45603 46461 45615 46464
rect 45557 46455 45615 46461
rect 38712 46396 40264 46424
rect 38712 46384 38718 46396
rect 41874 46384 41880 46436
rect 41932 46424 41938 46436
rect 43088 46424 43116 46455
rect 48038 46452 48044 46464
rect 48096 46452 48102 46504
rect 41932 46396 43116 46424
rect 41932 46384 41938 46396
rect 10410 46316 10416 46368
rect 10468 46356 10474 46368
rect 10689 46359 10747 46365
rect 10689 46356 10701 46359
rect 10468 46328 10701 46356
rect 10468 46316 10474 46328
rect 10689 46325 10701 46328
rect 10735 46325 10747 46359
rect 10689 46319 10747 46325
rect 22738 46316 22744 46368
rect 22796 46356 22802 46368
rect 29730 46356 29736 46368
rect 22796 46328 29736 46356
rect 22796 46316 22802 46328
rect 29730 46316 29736 46328
rect 29788 46316 29794 46368
rect 35526 46316 35532 46368
rect 35584 46356 35590 46368
rect 35805 46359 35863 46365
rect 35805 46356 35817 46359
rect 35584 46328 35817 46356
rect 35584 46316 35590 46328
rect 35805 46325 35817 46328
rect 35851 46325 35863 46359
rect 35805 46319 35863 46325
rect 45738 46316 45744 46368
rect 45796 46356 45802 46368
rect 47949 46359 48007 46365
rect 47949 46356 47961 46359
rect 45796 46328 47961 46356
rect 45796 46316 45802 46328
rect 47949 46325 47961 46328
rect 47995 46325 48007 46359
rect 47949 46319 48007 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 4890 46112 4896 46164
rect 4948 46152 4954 46164
rect 22738 46152 22744 46164
rect 4948 46124 22744 46152
rect 4948 46112 4954 46124
rect 22738 46112 22744 46124
rect 22796 46112 22802 46164
rect 22922 46152 22928 46164
rect 22883 46124 22928 46152
rect 22922 46112 22928 46124
rect 22980 46112 22986 46164
rect 26970 46152 26976 46164
rect 26931 46124 26976 46152
rect 26970 46112 26976 46124
rect 27028 46112 27034 46164
rect 29089 46155 29147 46161
rect 29089 46121 29101 46155
rect 29135 46152 29147 46155
rect 29638 46152 29644 46164
rect 29135 46124 29644 46152
rect 29135 46121 29147 46124
rect 29089 46115 29147 46121
rect 29638 46112 29644 46124
rect 29696 46112 29702 46164
rect 33226 46152 33232 46164
rect 33187 46124 33232 46152
rect 33226 46112 33232 46124
rect 33284 46112 33290 46164
rect 38013 46155 38071 46161
rect 38013 46121 38025 46155
rect 38059 46152 38071 46155
rect 39942 46152 39948 46164
rect 38059 46124 39948 46152
rect 38059 46121 38071 46124
rect 38013 46115 38071 46121
rect 39942 46112 39948 46124
rect 40000 46112 40006 46164
rect 44545 46155 44603 46161
rect 44545 46121 44557 46155
rect 44591 46152 44603 46155
rect 45554 46152 45560 46164
rect 44591 46124 45560 46152
rect 44591 46121 44603 46124
rect 44545 46115 44603 46121
rect 45554 46112 45560 46124
rect 45612 46112 45618 46164
rect 48038 46112 48044 46164
rect 48096 46152 48102 46164
rect 48133 46155 48191 46161
rect 48133 46152 48145 46155
rect 48096 46124 48145 46152
rect 48096 46112 48102 46124
rect 48133 46121 48145 46124
rect 48179 46121 48191 46155
rect 48133 46115 48191 46121
rect 14642 46044 14648 46096
rect 14700 46084 14706 46096
rect 16669 46087 16727 46093
rect 16669 46084 16681 46087
rect 14700 46056 16681 46084
rect 14700 46044 14706 46056
rect 16669 46053 16681 46056
rect 16715 46053 16727 46087
rect 41506 46084 41512 46096
rect 16669 46047 16727 46053
rect 22066 46056 41512 46084
rect 1762 46016 1768 46028
rect 1723 45988 1768 46016
rect 1762 45976 1768 45988
rect 1820 45976 1826 46028
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 4890 46016 4896 46028
rect 4851 45988 4896 46016
rect 4890 45976 4896 45988
rect 4948 45976 4954 46028
rect 5534 45976 5540 46028
rect 5592 46016 5598 46028
rect 5629 46019 5687 46025
rect 5629 46016 5641 46019
rect 5592 45988 5641 46016
rect 5592 45976 5598 45988
rect 5629 45985 5641 45988
rect 5675 45985 5687 46019
rect 5629 45979 5687 45985
rect 5810 45976 5816 46028
rect 5868 46016 5874 46028
rect 6089 46019 6147 46025
rect 6089 46016 6101 46019
rect 5868 45988 6101 46016
rect 5868 45976 5874 45988
rect 6089 45985 6101 45988
rect 6135 45985 6147 46019
rect 10410 46016 10416 46028
rect 10371 45988 10416 46016
rect 6089 45979 6147 45985
rect 10410 45976 10416 45988
rect 10468 45976 10474 46028
rect 10962 45976 10968 46028
rect 11020 46016 11026 46028
rect 11057 46019 11115 46025
rect 11057 46016 11069 46019
rect 11020 45988 11069 46016
rect 11020 45976 11026 45988
rect 11057 45985 11069 45988
rect 11103 45985 11115 46019
rect 11057 45979 11115 45985
rect 14277 46019 14335 46025
rect 14277 45985 14289 46019
rect 14323 46016 14335 46019
rect 14550 46016 14556 46028
rect 14323 45988 14556 46016
rect 14323 45985 14335 45988
rect 14277 45979 14335 45985
rect 14550 45976 14556 45988
rect 14608 45976 14614 46028
rect 14826 46016 14832 46028
rect 14787 45988 14832 46016
rect 14826 45976 14832 45988
rect 14884 45976 14890 46028
rect 1581 45951 1639 45957
rect 1581 45917 1593 45951
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 4341 45951 4399 45957
rect 4341 45917 4353 45951
rect 4387 45948 4399 45951
rect 4798 45948 4804 45960
rect 4387 45920 4804 45948
rect 4387 45917 4399 45920
rect 4341 45911 4399 45917
rect 1596 45880 1624 45911
rect 4798 45908 4804 45920
rect 4856 45908 4862 45960
rect 13081 45951 13139 45957
rect 13081 45917 13093 45951
rect 13127 45948 13139 45951
rect 13354 45948 13360 45960
rect 13127 45920 13360 45948
rect 13127 45917 13139 45920
rect 13081 45911 13139 45917
rect 13354 45908 13360 45920
rect 13412 45908 13418 45960
rect 13538 45948 13544 45960
rect 13499 45920 13544 45948
rect 13538 45908 13544 45920
rect 13596 45908 13602 45960
rect 16574 45948 16580 45960
rect 16487 45920 16580 45948
rect 16574 45908 16580 45920
rect 16632 45948 16638 45960
rect 22066 45948 22094 46056
rect 41506 46044 41512 46056
rect 41564 46044 41570 46096
rect 43993 46087 44051 46093
rect 43993 46053 44005 46087
rect 44039 46084 44051 46087
rect 45370 46084 45376 46096
rect 44039 46056 45376 46084
rect 44039 46053 44051 46056
rect 43993 46047 44051 46053
rect 45370 46044 45376 46056
rect 45428 46044 45434 46096
rect 47026 46044 47032 46096
rect 47084 46044 47090 46096
rect 25130 46016 25136 46028
rect 25091 45988 25136 46016
rect 25130 45976 25136 45988
rect 25188 45976 25194 46028
rect 29733 46019 29791 46025
rect 29733 45985 29745 46019
rect 29779 46016 29791 46019
rect 29914 46016 29920 46028
rect 29779 45988 29920 46016
rect 29779 45985 29791 45988
rect 29733 45979 29791 45985
rect 29914 45976 29920 45988
rect 29972 45976 29978 46028
rect 30282 45976 30288 46028
rect 30340 46016 30346 46028
rect 30377 46019 30435 46025
rect 30377 46016 30389 46019
rect 30340 45988 30389 46016
rect 30340 45976 30346 45988
rect 30377 45985 30389 45988
rect 30423 45985 30435 46019
rect 35526 46016 35532 46028
rect 35487 45988 35532 46016
rect 30377 45979 30435 45985
rect 35526 45976 35532 45988
rect 35584 45976 35590 46028
rect 36078 46016 36084 46028
rect 36039 45988 36084 46016
rect 36078 45976 36084 45988
rect 36136 45976 36142 46028
rect 40586 46016 40592 46028
rect 40547 45988 40592 46016
rect 40586 45976 40592 45988
rect 40644 45976 40650 46028
rect 45738 46016 45744 46028
rect 45699 45988 45744 46016
rect 45738 45976 45744 45988
rect 45796 45976 45802 46028
rect 47044 46016 47072 46044
rect 47121 46019 47179 46025
rect 47121 46016 47133 46019
rect 47044 45988 47133 46016
rect 47121 45985 47133 45988
rect 47167 45985 47179 46019
rect 47121 45979 47179 45985
rect 16632 45920 22094 45948
rect 22833 45951 22891 45957
rect 16632 45908 16638 45920
rect 22833 45917 22845 45951
rect 22879 45917 22891 45951
rect 22833 45911 22891 45917
rect 24029 45951 24087 45957
rect 24029 45917 24041 45951
rect 24075 45948 24087 45951
rect 24581 45951 24639 45957
rect 24581 45948 24593 45951
rect 24075 45920 24593 45948
rect 24075 45917 24087 45920
rect 24029 45911 24087 45917
rect 24581 45917 24593 45920
rect 24627 45917 24639 45951
rect 24581 45911 24639 45917
rect 26881 45951 26939 45957
rect 26881 45917 26893 45951
rect 26927 45948 26939 45951
rect 26970 45948 26976 45960
rect 26927 45920 26976 45948
rect 26927 45917 26939 45920
rect 26881 45911 26939 45917
rect 3050 45880 3056 45892
rect 1596 45852 3056 45880
rect 3050 45840 3056 45852
rect 3108 45840 3114 45892
rect 5813 45883 5871 45889
rect 5813 45849 5825 45883
rect 5859 45880 5871 45883
rect 6638 45880 6644 45892
rect 5859 45852 6644 45880
rect 5859 45849 5871 45852
rect 5813 45843 5871 45849
rect 6638 45840 6644 45852
rect 6696 45840 6702 45892
rect 10594 45880 10600 45892
rect 10555 45852 10600 45880
rect 10594 45840 10600 45852
rect 10652 45840 10658 45892
rect 13633 45883 13691 45889
rect 13633 45849 13645 45883
rect 13679 45880 13691 45883
rect 14461 45883 14519 45889
rect 14461 45880 14473 45883
rect 13679 45852 14473 45880
rect 13679 45849 13691 45852
rect 13633 45843 13691 45849
rect 14461 45849 14473 45852
rect 14507 45849 14519 45883
rect 14461 45843 14519 45849
rect 22848 45824 22876 45911
rect 26970 45908 26976 45920
rect 27028 45908 27034 45960
rect 28994 45948 29000 45960
rect 28955 45920 29000 45948
rect 28994 45908 29000 45920
rect 29052 45908 29058 45960
rect 33137 45951 33195 45957
rect 33137 45917 33149 45951
rect 33183 45917 33195 45951
rect 37918 45948 37924 45960
rect 37879 45920 37924 45948
rect 33137 45911 33195 45917
rect 24762 45880 24768 45892
rect 24723 45852 24768 45880
rect 24762 45840 24768 45852
rect 24820 45840 24826 45892
rect 29914 45880 29920 45892
rect 29875 45852 29920 45880
rect 29914 45840 29920 45852
rect 29972 45840 29978 45892
rect 22830 45812 22836 45824
rect 22743 45784 22836 45812
rect 22830 45772 22836 45784
rect 22888 45812 22894 45824
rect 33152 45812 33180 45911
rect 37918 45908 37924 45920
rect 37976 45908 37982 45960
rect 40126 45948 40132 45960
rect 40087 45920 40132 45948
rect 40126 45908 40132 45920
rect 40184 45908 40190 45960
rect 44453 45951 44511 45957
rect 44453 45917 44465 45951
rect 44499 45917 44511 45951
rect 48041 45951 48099 45957
rect 48041 45948 48053 45951
rect 44453 45911 44511 45917
rect 47596 45920 48053 45948
rect 35710 45880 35716 45892
rect 35671 45852 35716 45880
rect 35710 45840 35716 45852
rect 35768 45840 35774 45892
rect 40310 45880 40316 45892
rect 35866 45852 40172 45880
rect 40271 45852 40316 45880
rect 35866 45812 35894 45852
rect 22888 45784 35894 45812
rect 40144 45812 40172 45852
rect 40310 45840 40316 45852
rect 40368 45840 40374 45892
rect 44468 45812 44496 45911
rect 45922 45880 45928 45892
rect 45883 45852 45928 45880
rect 45922 45840 45928 45852
rect 45980 45840 45986 45892
rect 47596 45824 47624 45920
rect 48041 45917 48053 45920
rect 48087 45917 48099 45951
rect 48041 45911 48099 45917
rect 47578 45812 47584 45824
rect 40144 45784 47584 45812
rect 22888 45772 22894 45784
rect 47578 45772 47584 45784
rect 47636 45772 47642 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 6638 45608 6644 45620
rect 6599 45580 6644 45608
rect 6638 45568 6644 45580
rect 6696 45568 6702 45620
rect 10594 45608 10600 45620
rect 10555 45580 10600 45608
rect 10594 45568 10600 45580
rect 10652 45568 10658 45620
rect 13538 45568 13544 45620
rect 13596 45608 13602 45620
rect 24489 45611 24547 45617
rect 13596 45580 24440 45608
rect 13596 45568 13602 45580
rect 12434 45500 12440 45552
rect 12492 45540 12498 45552
rect 13081 45543 13139 45549
rect 12492 45512 12537 45540
rect 12492 45500 12498 45512
rect 13081 45509 13093 45543
rect 13127 45540 13139 45543
rect 13817 45543 13875 45549
rect 13817 45540 13829 45543
rect 13127 45512 13829 45540
rect 13127 45509 13139 45512
rect 13081 45503 13139 45509
rect 13817 45509 13829 45512
rect 13863 45509 13875 45543
rect 13817 45503 13875 45509
rect 4706 45472 4712 45484
rect 4667 45444 4712 45472
rect 4706 45432 4712 45444
rect 4764 45432 4770 45484
rect 4890 45432 4896 45484
rect 4948 45472 4954 45484
rect 6549 45475 6607 45481
rect 6549 45472 6561 45475
rect 4948 45444 6561 45472
rect 4948 45432 4954 45444
rect 6549 45441 6561 45444
rect 6595 45472 6607 45475
rect 6595 45444 10456 45472
rect 6595 45441 6607 45444
rect 6549 45435 6607 45441
rect 2225 45407 2283 45413
rect 2225 45373 2237 45407
rect 2271 45373 2283 45407
rect 2225 45367 2283 45373
rect 2409 45407 2467 45413
rect 2409 45373 2421 45407
rect 2455 45404 2467 45407
rect 2498 45404 2504 45416
rect 2455 45376 2504 45404
rect 2455 45373 2467 45376
rect 2409 45367 2467 45373
rect 2240 45336 2268 45367
rect 2498 45364 2504 45376
rect 2556 45364 2562 45416
rect 2958 45404 2964 45416
rect 2919 45376 2964 45404
rect 2958 45364 2964 45376
rect 3016 45364 3022 45416
rect 4982 45404 4988 45416
rect 4943 45376 4988 45404
rect 4982 45364 4988 45376
rect 5040 45404 5046 45416
rect 10318 45404 10324 45416
rect 5040 45376 10324 45404
rect 5040 45364 5046 45376
rect 10318 45364 10324 45376
rect 10376 45364 10382 45416
rect 2314 45336 2320 45348
rect 2240 45308 2320 45336
rect 2314 45296 2320 45308
rect 2372 45296 2378 45348
rect 10428 45336 10456 45444
rect 10502 45432 10508 45484
rect 10560 45472 10566 45484
rect 12342 45472 12348 45484
rect 10560 45444 10605 45472
rect 12303 45444 12348 45472
rect 10560 45432 10566 45444
rect 12342 45432 12348 45444
rect 12400 45432 12406 45484
rect 12986 45472 12992 45484
rect 12947 45444 12992 45472
rect 12986 45432 12992 45444
rect 13044 45432 13050 45484
rect 13354 45432 13360 45484
rect 13412 45472 13418 45484
rect 24412 45481 24440 45580
rect 24489 45577 24501 45611
rect 24535 45608 24547 45611
rect 24762 45608 24768 45620
rect 24535 45580 24768 45608
rect 24535 45577 24547 45580
rect 24489 45571 24547 45577
rect 24762 45568 24768 45580
rect 24820 45568 24826 45620
rect 24946 45568 24952 45620
rect 25004 45608 25010 45620
rect 25317 45611 25375 45617
rect 25317 45608 25329 45611
rect 25004 45580 25329 45608
rect 25004 45568 25010 45580
rect 25317 45577 25329 45580
rect 25363 45577 25375 45611
rect 25317 45571 25375 45577
rect 29825 45611 29883 45617
rect 29825 45577 29837 45611
rect 29871 45608 29883 45611
rect 29914 45608 29920 45620
rect 29871 45580 29920 45608
rect 29871 45577 29883 45580
rect 29825 45571 29883 45577
rect 29914 45568 29920 45580
rect 29972 45568 29978 45620
rect 35710 45608 35716 45620
rect 30024 45580 34560 45608
rect 35671 45580 35716 45608
rect 28994 45500 29000 45552
rect 29052 45540 29058 45552
rect 30024 45540 30052 45580
rect 29052 45512 30052 45540
rect 29052 45500 29058 45512
rect 13633 45475 13691 45481
rect 13633 45472 13645 45475
rect 13412 45444 13645 45472
rect 13412 45432 13418 45444
rect 13633 45441 13645 45444
rect 13679 45441 13691 45475
rect 13633 45435 13691 45441
rect 24397 45475 24455 45481
rect 24397 45441 24409 45475
rect 24443 45472 24455 45475
rect 25225 45475 25283 45481
rect 25225 45472 25237 45475
rect 24443 45444 25237 45472
rect 24443 45441 24455 45444
rect 24397 45435 24455 45441
rect 25225 45441 25237 45444
rect 25271 45472 25283 45475
rect 29012 45472 29040 45500
rect 29730 45472 29736 45484
rect 25271 45444 29040 45472
rect 29691 45444 29736 45472
rect 25271 45441 25283 45444
rect 25225 45435 25283 45441
rect 29730 45432 29736 45444
rect 29788 45432 29794 45484
rect 34532 45472 34560 45580
rect 35710 45568 35716 45580
rect 35768 45568 35774 45620
rect 36633 45543 36691 45549
rect 36633 45509 36645 45543
rect 36679 45540 36691 45543
rect 37642 45540 37648 45552
rect 36679 45512 37648 45540
rect 36679 45509 36691 45512
rect 36633 45503 36691 45509
rect 37642 45500 37648 45512
rect 37700 45500 37706 45552
rect 41601 45543 41659 45549
rect 41601 45509 41613 45543
rect 41647 45540 41659 45543
rect 42794 45540 42800 45552
rect 41647 45512 42800 45540
rect 41647 45509 41659 45512
rect 41601 45503 41659 45509
rect 42794 45500 42800 45512
rect 42852 45500 42858 45552
rect 45557 45543 45615 45549
rect 45557 45509 45569 45543
rect 45603 45540 45615 45543
rect 47854 45540 47860 45552
rect 45603 45512 47860 45540
rect 45603 45509 45615 45512
rect 45557 45503 45615 45509
rect 47854 45500 47860 45512
rect 47912 45500 47918 45552
rect 35618 45472 35624 45484
rect 34532 45444 35624 45472
rect 35618 45432 35624 45444
rect 35676 45432 35682 45484
rect 36538 45472 36544 45484
rect 36499 45444 36544 45472
rect 36538 45432 36544 45444
rect 36596 45472 36602 45484
rect 37918 45472 37924 45484
rect 36596 45444 37924 45472
rect 36596 45432 36602 45444
rect 37918 45432 37924 45444
rect 37976 45432 37982 45484
rect 40126 45432 40132 45484
rect 40184 45472 40190 45484
rect 40405 45475 40463 45481
rect 40405 45472 40417 45475
rect 40184 45444 40417 45472
rect 40184 45432 40190 45444
rect 40405 45441 40417 45444
rect 40451 45441 40463 45475
rect 41506 45472 41512 45484
rect 41467 45444 41512 45472
rect 40405 45435 40463 45441
rect 41506 45432 41512 45444
rect 41564 45432 41570 45484
rect 14182 45404 14188 45416
rect 14143 45376 14188 45404
rect 14182 45364 14188 45376
rect 14240 45364 14246 45416
rect 44913 45407 44971 45413
rect 44913 45373 44925 45407
rect 44959 45404 44971 45407
rect 45373 45407 45431 45413
rect 45373 45404 45385 45407
rect 44959 45376 45385 45404
rect 44959 45373 44971 45376
rect 44913 45367 44971 45373
rect 45373 45373 45385 45376
rect 45419 45373 45431 45407
rect 46842 45404 46848 45416
rect 46803 45376 46848 45404
rect 45373 45367 45431 45373
rect 46842 45364 46848 45376
rect 46900 45364 46906 45416
rect 26970 45336 26976 45348
rect 10428 45308 26976 45336
rect 26970 45296 26976 45308
rect 27028 45296 27034 45348
rect 1765 45271 1823 45277
rect 1765 45237 1777 45271
rect 1811 45268 1823 45271
rect 2222 45268 2228 45280
rect 1811 45240 2228 45268
rect 1811 45237 1823 45240
rect 1765 45231 1823 45237
rect 2222 45228 2228 45240
rect 2280 45228 2286 45280
rect 12342 45228 12348 45280
rect 12400 45268 12406 45280
rect 16574 45268 16580 45280
rect 12400 45240 16580 45268
rect 12400 45228 12406 45240
rect 16574 45228 16580 45240
rect 16632 45228 16638 45280
rect 46474 45228 46480 45280
rect 46532 45268 46538 45280
rect 47949 45271 48007 45277
rect 47949 45268 47961 45271
rect 46532 45240 47961 45268
rect 46532 45228 46538 45240
rect 47949 45237 47961 45240
rect 47995 45237 48007 45271
rect 47949 45231 48007 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 4433 45067 4491 45073
rect 4433 45033 4445 45067
rect 4479 45064 4491 45067
rect 4614 45064 4620 45076
rect 4479 45036 4620 45064
rect 4479 45033 4491 45036
rect 4433 45027 4491 45033
rect 4614 45024 4620 45036
rect 4672 45024 4678 45076
rect 40310 45064 40316 45076
rect 40271 45036 40316 45064
rect 40310 45024 40316 45036
rect 40368 45024 40374 45076
rect 45833 45067 45891 45073
rect 45833 45033 45845 45067
rect 45879 45064 45891 45067
rect 45922 45064 45928 45076
rect 45879 45036 45928 45064
rect 45879 45033 45891 45036
rect 45833 45027 45891 45033
rect 45922 45024 45928 45036
rect 45980 45024 45986 45076
rect 22830 44928 22836 44940
rect 3252 44900 22836 44928
rect 1762 44860 1768 44872
rect 1723 44832 1768 44860
rect 1762 44820 1768 44832
rect 1820 44820 1826 44872
rect 2593 44863 2651 44869
rect 2593 44829 2605 44863
rect 2639 44829 2651 44863
rect 2593 44823 2651 44829
rect 1857 44727 1915 44733
rect 1857 44693 1869 44727
rect 1903 44724 1915 44727
rect 2406 44724 2412 44736
rect 1903 44696 2412 44724
rect 1903 44693 1915 44696
rect 1857 44687 1915 44693
rect 2406 44684 2412 44696
rect 2464 44684 2470 44736
rect 2608 44724 2636 44823
rect 3252 44804 3280 44900
rect 22830 44888 22836 44900
rect 22888 44888 22894 44940
rect 46474 44928 46480 44940
rect 46435 44900 46480 44928
rect 46474 44888 46480 44900
rect 46532 44888 46538 44940
rect 48222 44928 48228 44940
rect 48183 44900 48228 44928
rect 48222 44888 48228 44900
rect 48280 44888 48286 44940
rect 4341 44863 4399 44869
rect 4341 44829 4353 44863
rect 4387 44860 4399 44863
rect 4890 44860 4896 44872
rect 4387 44832 4896 44860
rect 4387 44829 4399 44832
rect 4341 44823 4399 44829
rect 4890 44820 4896 44832
rect 4948 44820 4954 44872
rect 4985 44863 5043 44869
rect 4985 44829 4997 44863
rect 5031 44829 5043 44863
rect 40218 44860 40224 44872
rect 40179 44832 40224 44860
rect 4985 44823 5043 44829
rect 3234 44792 3240 44804
rect 3195 44764 3240 44792
rect 3234 44752 3240 44764
rect 3292 44752 3298 44804
rect 5000 44792 5028 44823
rect 40218 44820 40224 44832
rect 40276 44820 40282 44872
rect 45741 44863 45799 44869
rect 45741 44829 45753 44863
rect 45787 44829 45799 44863
rect 45741 44823 45799 44829
rect 4908 44764 5028 44792
rect 4522 44724 4528 44736
rect 2608 44696 4528 44724
rect 4522 44684 4528 44696
rect 4580 44724 4586 44736
rect 4706 44724 4712 44736
rect 4580 44696 4712 44724
rect 4580 44684 4586 44696
rect 4706 44684 4712 44696
rect 4764 44724 4770 44736
rect 4908 44724 4936 44764
rect 5718 44752 5724 44804
rect 5776 44792 5782 44804
rect 5813 44795 5871 44801
rect 5813 44792 5825 44795
rect 5776 44764 5825 44792
rect 5776 44752 5782 44764
rect 5813 44761 5825 44764
rect 5859 44792 5871 44795
rect 12342 44792 12348 44804
rect 5859 44764 12348 44792
rect 5859 44761 5871 44764
rect 5813 44755 5871 44761
rect 12342 44752 12348 44764
rect 12400 44752 12406 44804
rect 4764 44696 4936 44724
rect 45756 44724 45784 44823
rect 46658 44792 46664 44804
rect 46619 44764 46664 44792
rect 46658 44752 46664 44764
rect 46716 44752 46722 44804
rect 47670 44724 47676 44736
rect 45756 44696 47676 44724
rect 4764 44684 4770 44696
rect 47670 44684 47676 44696
rect 47728 44684 47734 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 1673 44523 1731 44529
rect 1673 44489 1685 44523
rect 1719 44520 1731 44523
rect 2498 44520 2504 44532
rect 1719 44492 2504 44520
rect 1719 44489 1731 44492
rect 1673 44483 1731 44489
rect 2498 44480 2504 44492
rect 2556 44480 2562 44532
rect 46477 44523 46535 44529
rect 46477 44489 46489 44523
rect 46523 44520 46535 44523
rect 46658 44520 46664 44532
rect 46523 44492 46664 44520
rect 46523 44489 46535 44492
rect 46477 44483 46535 44489
rect 46658 44480 46664 44492
rect 46716 44480 46722 44532
rect 2406 44452 2412 44464
rect 2367 44424 2412 44452
rect 2406 44412 2412 44424
rect 2464 44412 2470 44464
rect 7374 44452 7380 44464
rect 7287 44424 7380 44452
rect 7374 44412 7380 44424
rect 7432 44452 7438 44464
rect 12986 44452 12992 44464
rect 7432 44424 12992 44452
rect 7432 44412 7438 44424
rect 12986 44412 12992 44424
rect 13044 44412 13050 44464
rect 1581 44387 1639 44393
rect 1581 44353 1593 44387
rect 1627 44384 1639 44387
rect 2222 44384 2228 44396
rect 1627 44356 2084 44384
rect 2183 44356 2228 44384
rect 1627 44353 1639 44356
rect 1581 44347 1639 44353
rect 2056 44248 2084 44356
rect 2222 44344 2228 44356
rect 2280 44344 2286 44396
rect 4522 44384 4528 44396
rect 4483 44356 4528 44384
rect 4522 44344 4528 44356
rect 4580 44384 4586 44396
rect 6549 44387 6607 44393
rect 6549 44384 6561 44387
rect 4580 44356 6561 44384
rect 4580 44344 4586 44356
rect 6549 44353 6561 44356
rect 6595 44353 6607 44387
rect 6549 44347 6607 44353
rect 6886 44356 12434 44384
rect 2774 44316 2780 44328
rect 2735 44288 2780 44316
rect 2774 44276 2780 44288
rect 2832 44276 2838 44328
rect 5442 44316 5448 44328
rect 5403 44288 5448 44316
rect 5442 44276 5448 44288
rect 5500 44316 5506 44328
rect 6886 44316 6914 44356
rect 5500 44288 6914 44316
rect 12406 44316 12434 44356
rect 41506 44344 41512 44396
rect 41564 44384 41570 44396
rect 46385 44387 46443 44393
rect 46385 44384 46397 44387
rect 41564 44356 46397 44384
rect 41564 44344 41570 44356
rect 46385 44353 46397 44356
rect 46431 44384 46443 44387
rect 47762 44384 47768 44396
rect 46431 44356 47768 44384
rect 46431 44353 46443 44356
rect 46385 44347 46443 44353
rect 47762 44344 47768 44356
rect 47820 44344 47826 44396
rect 48314 44384 48320 44396
rect 48275 44356 48320 44384
rect 48314 44344 48320 44356
rect 48372 44344 48378 44396
rect 40218 44316 40224 44328
rect 12406 44288 40224 44316
rect 5500 44276 5506 44288
rect 40218 44276 40224 44288
rect 40276 44276 40282 44328
rect 3970 44248 3976 44260
rect 2056 44220 3976 44248
rect 3970 44208 3976 44220
rect 4028 44208 4034 44260
rect 47210 44180 47216 44192
rect 47171 44152 47216 44180
rect 47210 44140 47216 44152
rect 47268 44140 47274 44192
rect 47302 44140 47308 44192
rect 47360 44180 47366 44192
rect 48133 44183 48191 44189
rect 48133 44180 48145 44183
rect 47360 44152 48145 44180
rect 47360 44140 47366 44152
rect 48133 44149 48145 44152
rect 48179 44149 48191 44183
rect 48133 44143 48191 44149
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 4062 43976 4068 43988
rect 4023 43948 4068 43976
rect 4062 43936 4068 43948
rect 4120 43936 4126 43988
rect 2774 43840 2780 43852
rect 2735 43812 2780 43840
rect 2774 43800 2780 43812
rect 2832 43800 2838 43852
rect 4982 43840 4988 43852
rect 3988 43812 4988 43840
rect 3988 43784 4016 43812
rect 4982 43800 4988 43812
rect 5040 43800 5046 43852
rect 5534 43840 5540 43852
rect 5495 43812 5540 43840
rect 5534 43800 5540 43812
rect 5592 43800 5598 43852
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 47210 43840 47216 43852
rect 46523 43812 47216 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 47210 43800 47216 43812
rect 47268 43800 47274 43852
rect 48130 43840 48136 43852
rect 48091 43812 48136 43840
rect 48130 43800 48136 43812
rect 48188 43800 48194 43852
rect 1578 43772 1584 43784
rect 1539 43744 1584 43772
rect 1578 43732 1584 43744
rect 1636 43732 1642 43784
rect 3970 43772 3976 43784
rect 3931 43744 3976 43772
rect 3970 43732 3976 43744
rect 4028 43732 4034 43784
rect 4706 43732 4712 43784
rect 4764 43772 4770 43784
rect 5077 43775 5135 43781
rect 5077 43772 5089 43775
rect 4764 43744 5089 43772
rect 4764 43732 4770 43744
rect 5077 43741 5089 43744
rect 5123 43741 5135 43775
rect 5077 43735 5135 43741
rect 27065 43775 27123 43781
rect 27065 43741 27077 43775
rect 27111 43741 27123 43775
rect 27065 43735 27123 43741
rect 27157 43775 27215 43781
rect 27157 43741 27169 43775
rect 27203 43772 27215 43775
rect 27798 43772 27804 43784
rect 27203 43744 27804 43772
rect 27203 43741 27215 43744
rect 27157 43735 27215 43741
rect 1765 43707 1823 43713
rect 1765 43673 1777 43707
rect 1811 43704 1823 43707
rect 2590 43704 2596 43716
rect 1811 43676 2596 43704
rect 1811 43673 1823 43676
rect 1765 43667 1823 43673
rect 2590 43664 2596 43676
rect 2648 43664 2654 43716
rect 5534 43664 5540 43716
rect 5592 43704 5598 43716
rect 13538 43704 13544 43716
rect 5592 43676 13544 43704
rect 5592 43664 5598 43676
rect 13538 43664 13544 43676
rect 13596 43664 13602 43716
rect 27080 43704 27108 43735
rect 27798 43732 27804 43744
rect 27856 43732 27862 43784
rect 27430 43704 27436 43716
rect 27080 43676 27436 43704
rect 27430 43664 27436 43676
rect 27488 43664 27494 43716
rect 46661 43707 46719 43713
rect 46661 43673 46673 43707
rect 46707 43704 46719 43707
rect 47118 43704 47124 43716
rect 46707 43676 47124 43704
rect 46707 43673 46719 43676
rect 46661 43667 46719 43673
rect 47118 43664 47124 43676
rect 47176 43664 47182 43716
rect 27338 43636 27344 43648
rect 27299 43608 27344 43636
rect 27338 43596 27344 43608
rect 27396 43596 27402 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 2590 43432 2596 43444
rect 2551 43404 2596 43432
rect 2590 43392 2596 43404
rect 2648 43392 2654 43444
rect 4614 43392 4620 43444
rect 4672 43432 4678 43444
rect 47118 43432 47124 43444
rect 4672 43404 45554 43432
rect 47079 43404 47124 43432
rect 4672 43392 4678 43404
rect 7834 43324 7840 43376
rect 7892 43364 7898 43376
rect 22281 43367 22339 43373
rect 22281 43364 22293 43367
rect 7892 43336 22293 43364
rect 7892 43324 7898 43336
rect 22281 43333 22293 43336
rect 22327 43364 22339 43367
rect 22370 43364 22376 43376
rect 22327 43336 22376 43364
rect 22327 43333 22339 43336
rect 22281 43327 22339 43333
rect 22370 43324 22376 43336
rect 22428 43324 22434 43376
rect 22480 43336 23704 43364
rect 1578 43256 1584 43308
rect 1636 43296 1642 43308
rect 2041 43299 2099 43305
rect 2041 43296 2053 43299
rect 1636 43268 2053 43296
rect 1636 43256 1642 43268
rect 2041 43265 2053 43268
rect 2087 43265 2099 43299
rect 2041 43259 2099 43265
rect 2501 43299 2559 43305
rect 2501 43265 2513 43299
rect 2547 43265 2559 43299
rect 2501 43259 2559 43265
rect 3881 43299 3939 43305
rect 3881 43265 3893 43299
rect 3927 43296 3939 43299
rect 4706 43296 4712 43308
rect 3927 43268 4712 43296
rect 3927 43265 3939 43268
rect 3881 43259 3939 43265
rect 1946 43188 1952 43240
rect 2004 43228 2010 43240
rect 2516 43228 2544 43259
rect 4706 43256 4712 43268
rect 4764 43256 4770 43308
rect 9122 43256 9128 43308
rect 9180 43296 9186 43308
rect 9180 43268 12434 43296
rect 9180 43256 9186 43268
rect 4614 43228 4620 43240
rect 2004 43200 2544 43228
rect 4575 43200 4620 43228
rect 2004 43188 2010 43200
rect 4614 43188 4620 43200
rect 4672 43188 4678 43240
rect 12406 43228 12434 43268
rect 22480 43228 22508 43336
rect 22554 43256 22560 43308
rect 22612 43294 22618 43308
rect 23676 43305 23704 43336
rect 29730 43324 29736 43376
rect 29788 43364 29794 43376
rect 29788 43336 36216 43364
rect 29788 43324 29794 43336
rect 22833 43299 22891 43305
rect 22833 43296 22845 43299
rect 22664 43294 22845 43296
rect 22612 43268 22845 43294
rect 22612 43266 22692 43268
rect 22612 43256 22618 43266
rect 22833 43265 22845 43268
rect 22879 43265 22891 43299
rect 22833 43259 22891 43265
rect 23661 43299 23719 43305
rect 23661 43265 23673 43299
rect 23707 43296 23719 43299
rect 24121 43299 24179 43305
rect 24121 43296 24133 43299
rect 23707 43268 24133 43296
rect 23707 43265 23719 43268
rect 23661 43259 23719 43265
rect 24121 43265 24133 43268
rect 24167 43265 24179 43299
rect 27338 43296 27344 43308
rect 27299 43268 27344 43296
rect 24121 43259 24179 43265
rect 27338 43256 27344 43268
rect 27396 43256 27402 43308
rect 28445 43299 28503 43305
rect 28445 43265 28457 43299
rect 28491 43296 28503 43299
rect 28534 43296 28540 43308
rect 28491 43268 28540 43296
rect 28491 43265 28503 43268
rect 28445 43259 28503 43265
rect 28534 43256 28540 43268
rect 28592 43256 28598 43308
rect 28712 43299 28770 43305
rect 28712 43265 28724 43299
rect 28758 43296 28770 43299
rect 28994 43296 29000 43308
rect 28758 43268 29000 43296
rect 28758 43265 28770 43268
rect 28712 43259 28770 43265
rect 28994 43256 29000 43268
rect 29052 43256 29058 43308
rect 30466 43296 30472 43308
rect 30427 43268 30472 43296
rect 30466 43256 30472 43268
rect 30524 43256 30530 43308
rect 35897 43299 35955 43305
rect 35897 43265 35909 43299
rect 35943 43296 35955 43299
rect 36078 43296 36084 43308
rect 35943 43268 36084 43296
rect 35943 43265 35955 43268
rect 35897 43259 35955 43265
rect 36078 43256 36084 43268
rect 36136 43256 36142 43308
rect 12406 43200 22508 43228
rect 22649 43231 22707 43237
rect 22649 43197 22661 43231
rect 22695 43228 22707 43231
rect 23845 43231 23903 43237
rect 23845 43228 23857 43231
rect 22695 43200 23857 43228
rect 22695 43197 22707 43200
rect 22649 43191 22707 43197
rect 23845 43197 23857 43200
rect 23891 43228 23903 43231
rect 27430 43228 27436 43240
rect 23891 43200 27436 43228
rect 23891 43197 23903 43200
rect 23845 43191 23903 43197
rect 27430 43188 27436 43200
rect 27488 43188 27494 43240
rect 36188 43228 36216 43336
rect 45526 43296 45554 43404
rect 47118 43392 47124 43404
rect 47176 43392 47182 43444
rect 47026 43296 47032 43308
rect 45526 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 47486 43256 47492 43308
rect 47544 43296 47550 43308
rect 47765 43299 47823 43305
rect 47765 43296 47777 43299
rect 47544 43268 47777 43296
rect 47544 43256 47550 43268
rect 47765 43265 47777 43268
rect 47811 43265 47823 43299
rect 47765 43259 47823 43265
rect 47504 43228 47532 43256
rect 36188 43200 47532 43228
rect 23017 43163 23075 43169
rect 23017 43129 23029 43163
rect 23063 43160 23075 43163
rect 23658 43160 23664 43172
rect 23063 43132 23664 43160
rect 23063 43129 23075 43132
rect 23017 43123 23075 43129
rect 23658 43120 23664 43132
rect 23716 43120 23722 43172
rect 23477 43095 23535 43101
rect 23477 43061 23489 43095
rect 23523 43092 23535 43095
rect 23566 43092 23572 43104
rect 23523 43064 23572 43092
rect 23523 43061 23535 43064
rect 23477 43055 23535 43061
rect 23566 43052 23572 43064
rect 23624 43052 23630 43104
rect 27157 43095 27215 43101
rect 27157 43061 27169 43095
rect 27203 43092 27215 43095
rect 27246 43092 27252 43104
rect 27203 43064 27252 43092
rect 27203 43061 27215 43064
rect 27157 43055 27215 43061
rect 27246 43052 27252 43064
rect 27304 43052 27310 43104
rect 29822 43092 29828 43104
rect 29783 43064 29828 43092
rect 29822 43052 29828 43064
rect 29880 43052 29886 43104
rect 30282 43092 30288 43104
rect 30243 43064 30288 43092
rect 30282 43052 30288 43064
rect 30340 43052 30346 43104
rect 35713 43095 35771 43101
rect 35713 43061 35725 43095
rect 35759 43092 35771 43095
rect 35894 43092 35900 43104
rect 35759 43064 35900 43092
rect 35759 43061 35771 43064
rect 35713 43055 35771 43061
rect 35894 43052 35900 43064
rect 35952 43052 35958 43104
rect 47854 43092 47860 43104
rect 47815 43064 47860 43092
rect 47854 43052 47860 43064
rect 47912 43052 47918 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 2314 42712 2320 42764
rect 2372 42752 2378 42764
rect 2409 42755 2467 42761
rect 2409 42752 2421 42755
rect 2372 42724 2421 42752
rect 2372 42712 2378 42724
rect 2409 42721 2421 42724
rect 2455 42721 2467 42755
rect 3050 42752 3056 42764
rect 3011 42724 3056 42752
rect 2409 42715 2467 42721
rect 3050 42712 3056 42724
rect 3108 42712 3114 42764
rect 4706 42752 4712 42764
rect 4667 42724 4712 42752
rect 4706 42712 4712 42724
rect 4764 42712 4770 42764
rect 28074 42712 28080 42764
rect 28132 42752 28138 42764
rect 28534 42752 28540 42764
rect 28132 42724 28540 42752
rect 28132 42712 28138 42724
rect 28534 42712 28540 42724
rect 28592 42752 28598 42764
rect 29733 42755 29791 42761
rect 29733 42752 29745 42755
rect 28592 42724 29745 42752
rect 28592 42712 28598 42724
rect 29733 42721 29745 42724
rect 29779 42721 29791 42755
rect 29733 42715 29791 42721
rect 46661 42755 46719 42761
rect 46661 42721 46673 42755
rect 46707 42752 46719 42755
rect 47854 42752 47860 42764
rect 46707 42724 47860 42752
rect 46707 42721 46719 42724
rect 46661 42715 46719 42721
rect 47854 42712 47860 42724
rect 47912 42712 47918 42764
rect 48222 42752 48228 42764
rect 48183 42724 48228 42752
rect 48222 42712 48228 42724
rect 48280 42712 48286 42764
rect 1765 42687 1823 42693
rect 1765 42653 1777 42687
rect 1811 42684 1823 42687
rect 2866 42684 2872 42696
rect 1811 42656 2872 42684
rect 1811 42653 1823 42656
rect 1765 42647 1823 42653
rect 2866 42644 2872 42656
rect 2924 42644 2930 42696
rect 4433 42687 4491 42693
rect 4433 42653 4445 42687
rect 4479 42684 4491 42687
rect 4798 42684 4804 42696
rect 4479 42656 4804 42684
rect 4479 42653 4491 42656
rect 4433 42647 4491 42653
rect 4798 42644 4804 42656
rect 4856 42644 4862 42696
rect 23658 42684 23664 42696
rect 23619 42656 23664 42684
rect 23658 42644 23664 42656
rect 23716 42644 23722 42696
rect 27525 42687 27583 42693
rect 27525 42653 27537 42687
rect 27571 42653 27583 42687
rect 28442 42684 28448 42696
rect 28403 42656 28448 42684
rect 27525 42647 27583 42653
rect 27540 42616 27568 42647
rect 28442 42644 28448 42656
rect 28500 42644 28506 42696
rect 28629 42687 28687 42693
rect 28629 42653 28641 42687
rect 28675 42684 28687 42687
rect 28718 42684 28724 42696
rect 28675 42656 28724 42684
rect 28675 42653 28687 42656
rect 28629 42647 28687 42653
rect 28718 42644 28724 42656
rect 28776 42644 28782 42696
rect 30000 42687 30058 42693
rect 30000 42653 30012 42687
rect 30046 42684 30058 42687
rect 30282 42684 30288 42696
rect 30046 42656 30288 42684
rect 30046 42653 30058 42656
rect 30000 42647 30058 42653
rect 30282 42644 30288 42656
rect 30340 42644 30346 42696
rect 31573 42687 31631 42693
rect 31573 42653 31585 42687
rect 31619 42684 31631 42687
rect 32122 42684 32128 42696
rect 31619 42656 32128 42684
rect 31619 42653 31631 42656
rect 31573 42647 31631 42653
rect 32122 42644 32128 42656
rect 32180 42684 32186 42696
rect 35069 42687 35127 42693
rect 32180 42656 33916 42684
rect 32180 42644 32186 42656
rect 33888 42628 33916 42656
rect 35069 42653 35081 42687
rect 35115 42684 35127 42687
rect 35342 42684 35348 42696
rect 35115 42656 35348 42684
rect 35115 42653 35127 42656
rect 35069 42647 35127 42653
rect 35342 42644 35348 42656
rect 35400 42644 35406 42696
rect 35805 42687 35863 42693
rect 35805 42653 35817 42687
rect 35851 42653 35863 42687
rect 35805 42647 35863 42653
rect 28902 42616 28908 42628
rect 27540 42588 28908 42616
rect 28902 42576 28908 42588
rect 28960 42576 28966 42628
rect 31840 42619 31898 42625
rect 31840 42585 31852 42619
rect 31886 42616 31898 42619
rect 32858 42616 32864 42628
rect 31886 42588 32864 42616
rect 31886 42585 31898 42588
rect 31840 42579 31898 42585
rect 32858 42576 32864 42588
rect 32916 42576 32922 42628
rect 33870 42576 33876 42628
rect 33928 42616 33934 42628
rect 35820 42616 35848 42647
rect 35894 42644 35900 42696
rect 35952 42684 35958 42696
rect 36061 42687 36119 42693
rect 36061 42684 36073 42687
rect 35952 42656 36073 42684
rect 35952 42644 35958 42656
rect 36061 42653 36073 42656
rect 36107 42653 36119 42687
rect 36061 42647 36119 42653
rect 46017 42687 46075 42693
rect 46017 42653 46029 42687
rect 46063 42684 46075 42687
rect 46477 42687 46535 42693
rect 46477 42684 46489 42687
rect 46063 42656 46489 42684
rect 46063 42653 46075 42656
rect 46017 42647 46075 42653
rect 46477 42653 46489 42656
rect 46523 42653 46535 42687
rect 46477 42647 46535 42653
rect 33928 42588 35848 42616
rect 33928 42576 33934 42588
rect 1581 42551 1639 42557
rect 1581 42517 1593 42551
rect 1627 42548 1639 42551
rect 2682 42548 2688 42560
rect 1627 42520 2688 42548
rect 1627 42517 1639 42520
rect 1581 42511 1639 42517
rect 2682 42508 2688 42520
rect 2740 42508 2746 42560
rect 23474 42548 23480 42560
rect 23435 42520 23480 42548
rect 23474 42508 23480 42520
rect 23532 42508 23538 42560
rect 27338 42548 27344 42560
rect 27299 42520 27344 42548
rect 27338 42508 27344 42520
rect 27396 42508 27402 42560
rect 28813 42551 28871 42557
rect 28813 42517 28825 42551
rect 28859 42548 28871 42551
rect 29178 42548 29184 42560
rect 28859 42520 29184 42548
rect 28859 42517 28871 42520
rect 28813 42511 28871 42517
rect 29178 42508 29184 42520
rect 29236 42508 29242 42560
rect 31110 42548 31116 42560
rect 31071 42520 31116 42548
rect 31110 42508 31116 42520
rect 31168 42508 31174 42560
rect 32398 42508 32404 42560
rect 32456 42548 32462 42560
rect 32953 42551 33011 42557
rect 32953 42548 32965 42551
rect 32456 42520 32965 42548
rect 32456 42508 32462 42520
rect 32953 42517 32965 42520
rect 32999 42517 33011 42551
rect 34882 42548 34888 42560
rect 34843 42520 34888 42548
rect 32953 42511 33011 42517
rect 34882 42508 34888 42520
rect 34940 42508 34946 42560
rect 37182 42548 37188 42560
rect 37143 42520 37188 42548
rect 37182 42508 37188 42520
rect 37240 42508 37246 42560
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 22066 42316 31754 42344
rect 4706 42236 4712 42288
rect 4764 42276 4770 42288
rect 22066 42276 22094 42316
rect 4764 42248 22094 42276
rect 4764 42236 4770 42248
rect 23474 42236 23480 42288
rect 23532 42276 23538 42288
rect 24458 42279 24516 42285
rect 24458 42276 24470 42279
rect 23532 42248 24470 42276
rect 23532 42236 23538 42248
rect 24458 42245 24470 42248
rect 24504 42245 24516 42279
rect 28074 42276 28080 42288
rect 24458 42239 24516 42245
rect 27172 42248 28080 42276
rect 23566 42208 23572 42220
rect 23527 42180 23572 42208
rect 23566 42168 23572 42180
rect 23624 42168 23630 42220
rect 24213 42211 24271 42217
rect 24213 42177 24225 42211
rect 24259 42208 24271 42211
rect 24302 42208 24308 42220
rect 24259 42180 24308 42208
rect 24259 42177 24271 42180
rect 24213 42171 24271 42177
rect 24302 42168 24308 42180
rect 24360 42168 24366 42220
rect 27172 42217 27200 42248
rect 28074 42236 28080 42248
rect 28132 42236 28138 42288
rect 28718 42236 28724 42288
rect 28776 42276 28782 42288
rect 30101 42279 30159 42285
rect 28776 42248 29960 42276
rect 28776 42236 28782 42248
rect 27157 42211 27215 42217
rect 27157 42177 27169 42211
rect 27203 42177 27215 42211
rect 27157 42171 27215 42177
rect 27246 42168 27252 42220
rect 27304 42208 27310 42220
rect 27413 42211 27471 42217
rect 27413 42208 27425 42211
rect 27304 42180 27425 42208
rect 27304 42168 27310 42180
rect 27413 42177 27425 42180
rect 27459 42177 27471 42211
rect 29178 42208 29184 42220
rect 29139 42180 29184 42208
rect 27413 42171 27471 42177
rect 29178 42168 29184 42180
rect 29236 42168 29242 42220
rect 29822 42208 29828 42220
rect 29783 42180 29828 42208
rect 29822 42168 29828 42180
rect 29880 42168 29886 42220
rect 29932 42217 29960 42248
rect 30101 42245 30113 42279
rect 30147 42276 30159 42279
rect 30466 42276 30472 42288
rect 30147 42248 30472 42276
rect 30147 42245 30159 42248
rect 30101 42239 30159 42245
rect 30466 42236 30472 42248
rect 30524 42236 30530 42288
rect 31726 42276 31754 42316
rect 32858 42304 32864 42356
rect 32916 42344 32922 42356
rect 32953 42347 33011 42353
rect 32953 42344 32965 42347
rect 32916 42316 32965 42344
rect 32916 42304 32922 42316
rect 32953 42313 32965 42316
rect 32999 42313 33011 42347
rect 36078 42344 36084 42356
rect 36039 42316 36084 42344
rect 32953 42307 33011 42313
rect 36078 42304 36084 42316
rect 36136 42304 36142 42356
rect 36538 42276 36544 42288
rect 30944 42248 31248 42276
rect 31726 42248 36544 42276
rect 29917 42211 29975 42217
rect 29917 42177 29929 42211
rect 29963 42208 29975 42211
rect 30944 42208 30972 42248
rect 31110 42208 31116 42220
rect 29963 42180 30972 42208
rect 31071 42180 31116 42208
rect 29963 42177 29975 42180
rect 29917 42171 29975 42177
rect 31110 42168 31116 42180
rect 31168 42168 31174 42220
rect 31220 42217 31248 42248
rect 36538 42236 36544 42248
rect 36596 42236 36602 42288
rect 37829 42279 37887 42285
rect 37829 42276 37841 42279
rect 36924 42248 37841 42276
rect 31205 42211 31263 42217
rect 31205 42177 31217 42211
rect 31251 42177 31263 42211
rect 32490 42208 32496 42220
rect 32451 42180 32496 42208
rect 31205 42171 31263 42177
rect 29840 42140 29868 42168
rect 30558 42140 30564 42152
rect 29840 42112 30564 42140
rect 30558 42100 30564 42112
rect 30616 42100 30622 42152
rect 28994 42072 29000 42084
rect 28955 42044 29000 42072
rect 28994 42032 29000 42044
rect 29052 42032 29058 42084
rect 31220 42072 31248 42171
rect 32490 42168 32496 42180
rect 32548 42168 32554 42220
rect 33137 42211 33195 42217
rect 33137 42177 33149 42211
rect 33183 42177 33195 42211
rect 33870 42208 33876 42220
rect 33831 42180 33876 42208
rect 33137 42171 33195 42177
rect 31389 42143 31447 42149
rect 31389 42109 31401 42143
rect 31435 42140 31447 42143
rect 33152 42140 33180 42171
rect 33870 42168 33876 42180
rect 33928 42168 33934 42220
rect 34140 42211 34198 42217
rect 34140 42177 34152 42211
rect 34186 42208 34198 42211
rect 34882 42208 34888 42220
rect 34186 42180 34888 42208
rect 34186 42177 34198 42180
rect 34140 42171 34198 42177
rect 34882 42168 34888 42180
rect 34940 42168 34946 42220
rect 35894 42168 35900 42220
rect 35952 42208 35958 42220
rect 36924 42217 36952 42248
rect 37829 42245 37841 42248
rect 37875 42245 37887 42279
rect 47302 42276 47308 42288
rect 37829 42239 37887 42245
rect 40052 42248 47308 42276
rect 36909 42211 36967 42217
rect 35952 42180 35997 42208
rect 35952 42168 35958 42180
rect 36909 42177 36921 42211
rect 36955 42177 36967 42211
rect 37642 42208 37648 42220
rect 37603 42180 37648 42208
rect 36909 42171 36967 42177
rect 37642 42168 37648 42180
rect 37700 42168 37706 42220
rect 38473 42211 38531 42217
rect 38473 42177 38485 42211
rect 38519 42208 38531 42211
rect 38562 42208 38568 42220
rect 38519 42180 38568 42208
rect 38519 42177 38531 42180
rect 38473 42171 38531 42177
rect 38562 42168 38568 42180
rect 38620 42168 38626 42220
rect 40052 42217 40080 42248
rect 47302 42236 47308 42248
rect 47360 42236 47366 42288
rect 40037 42211 40095 42217
rect 40037 42177 40049 42211
rect 40083 42177 40095 42211
rect 40037 42171 40095 42177
rect 42880 42211 42938 42217
rect 42880 42177 42892 42211
rect 42926 42208 42938 42211
rect 43438 42208 43444 42220
rect 42926 42180 43444 42208
rect 42926 42177 42938 42180
rect 42880 42171 42938 42177
rect 43438 42168 43444 42180
rect 43496 42168 43502 42220
rect 47762 42208 47768 42220
rect 47723 42180 47768 42208
rect 47762 42168 47768 42180
rect 47820 42168 47826 42220
rect 35713 42143 35771 42149
rect 35713 42140 35725 42143
rect 31435 42112 33180 42140
rect 35544 42112 35725 42140
rect 31435 42109 31447 42112
rect 31389 42103 31447 42109
rect 33134 42072 33140 42084
rect 31220 42044 33140 42072
rect 33134 42032 33140 42044
rect 33192 42032 33198 42084
rect 35544 42016 35572 42112
rect 35713 42109 35725 42112
rect 35759 42109 35771 42143
rect 35713 42103 35771 42109
rect 37182 42100 37188 42152
rect 37240 42140 37246 42152
rect 37461 42143 37519 42149
rect 37461 42140 37473 42143
rect 37240 42112 37473 42140
rect 37240 42100 37246 42112
rect 37461 42109 37473 42112
rect 37507 42109 37519 42143
rect 37461 42103 37519 42109
rect 38746 42100 38752 42152
rect 38804 42140 38810 42152
rect 39853 42143 39911 42149
rect 39853 42140 39865 42143
rect 38804 42112 39865 42140
rect 38804 42100 38810 42112
rect 39853 42109 39865 42112
rect 39899 42109 39911 42143
rect 42610 42140 42616 42152
rect 42571 42112 42616 42140
rect 39853 42103 39911 42109
rect 42610 42100 42616 42112
rect 42668 42100 42674 42152
rect 23382 42004 23388 42016
rect 23343 41976 23388 42004
rect 23382 41964 23388 41976
rect 23440 41964 23446 42016
rect 25593 42007 25651 42013
rect 25593 41973 25605 42007
rect 25639 42004 25651 42007
rect 27890 42004 27896 42016
rect 25639 41976 27896 42004
rect 25639 41973 25651 41976
rect 25593 41967 25651 41973
rect 27890 41964 27896 41976
rect 27948 41964 27954 42016
rect 28534 42004 28540 42016
rect 28495 41976 28540 42004
rect 28534 41964 28540 41976
rect 28592 41964 28598 42016
rect 32306 42004 32312 42016
rect 32267 41976 32312 42004
rect 32306 41964 32312 41976
rect 32364 41964 32370 42016
rect 35253 42007 35311 42013
rect 35253 41973 35265 42007
rect 35299 42004 35311 42007
rect 35526 42004 35532 42016
rect 35299 41976 35532 42004
rect 35299 41973 35311 41976
rect 35253 41967 35311 41973
rect 35526 41964 35532 41976
rect 35584 41964 35590 42016
rect 36722 42004 36728 42016
rect 36683 41976 36728 42004
rect 36722 41964 36728 41976
rect 36780 41964 36786 42016
rect 38286 42004 38292 42016
rect 38247 41976 38292 42004
rect 38286 41964 38292 41976
rect 38344 41964 38350 42016
rect 40218 42004 40224 42016
rect 40179 41976 40224 42004
rect 40218 41964 40224 41976
rect 40276 41964 40282 42016
rect 43990 42004 43996 42016
rect 43951 41976 43996 42004
rect 43990 41964 43996 41976
rect 44048 41964 44054 42016
rect 46474 41964 46480 42016
rect 46532 42004 46538 42016
rect 47213 42007 47271 42013
rect 47213 42004 47225 42007
rect 46532 41976 47225 42004
rect 46532 41964 46538 41976
rect 47213 41973 47225 41976
rect 47259 41973 47271 42007
rect 47854 42004 47860 42016
rect 47815 41976 47860 42004
rect 47213 41967 47271 41973
rect 47854 41964 47860 41976
rect 47912 41964 47918 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 25961 41803 26019 41809
rect 25961 41769 25973 41803
rect 26007 41800 26019 41803
rect 28077 41803 28135 41809
rect 26007 41772 28028 41800
rect 26007 41769 26019 41772
rect 25961 41763 26019 41769
rect 28000 41732 28028 41772
rect 28077 41769 28089 41803
rect 28123 41800 28135 41803
rect 28442 41800 28448 41812
rect 28123 41772 28448 41800
rect 28123 41769 28135 41772
rect 28077 41763 28135 41769
rect 28442 41760 28448 41772
rect 28500 41800 28506 41812
rect 28626 41800 28632 41812
rect 28500 41772 28632 41800
rect 28500 41760 28506 41772
rect 28626 41760 28632 41772
rect 28684 41760 28690 41812
rect 28902 41800 28908 41812
rect 28863 41772 28908 41800
rect 28902 41760 28908 41772
rect 28960 41760 28966 41812
rect 35253 41803 35311 41809
rect 35253 41769 35265 41803
rect 35299 41800 35311 41803
rect 35342 41800 35348 41812
rect 35299 41772 35348 41800
rect 35299 41769 35311 41772
rect 35253 41763 35311 41769
rect 35342 41760 35348 41772
rect 35400 41760 35406 41812
rect 35894 41800 35900 41812
rect 35866 41760 35900 41800
rect 35952 41800 35958 41812
rect 37642 41800 37648 41812
rect 35952 41772 37648 41800
rect 35952 41760 35958 41772
rect 37642 41760 37648 41772
rect 37700 41760 37706 41812
rect 38562 41800 38568 41812
rect 38523 41772 38568 41800
rect 38562 41760 38568 41772
rect 38620 41760 38626 41812
rect 43438 41760 43444 41812
rect 43496 41800 43502 41812
rect 43533 41803 43591 41809
rect 43533 41800 43545 41803
rect 43496 41772 43545 41800
rect 43496 41760 43502 41772
rect 43533 41769 43545 41772
rect 43579 41769 43591 41803
rect 43533 41763 43591 41769
rect 30561 41735 30619 41741
rect 28000 41704 28994 41732
rect 28966 41664 28994 41704
rect 30561 41701 30573 41735
rect 30607 41732 30619 41735
rect 31110 41732 31116 41744
rect 30607 41704 31116 41732
rect 30607 41701 30619 41704
rect 30561 41695 30619 41701
rect 31110 41692 31116 41704
rect 31168 41692 31174 41744
rect 31478 41664 31484 41676
rect 28966 41636 31484 41664
rect 31478 41624 31484 41636
rect 31536 41624 31542 41676
rect 2038 41556 2044 41608
rect 2096 41596 2102 41608
rect 2317 41599 2375 41605
rect 2317 41596 2329 41599
rect 2096 41568 2329 41596
rect 2096 41556 2102 41568
rect 2317 41565 2329 41568
rect 2363 41565 2375 41599
rect 2317 41559 2375 41565
rect 24302 41556 24308 41608
rect 24360 41596 24366 41608
rect 24581 41599 24639 41605
rect 24581 41596 24593 41599
rect 24360 41568 24593 41596
rect 24360 41556 24366 41568
rect 24581 41565 24593 41568
rect 24627 41596 24639 41599
rect 26697 41599 26755 41605
rect 26697 41596 26709 41599
rect 24627 41568 26709 41596
rect 24627 41565 24639 41568
rect 24581 41559 24639 41565
rect 26697 41565 26709 41568
rect 26743 41596 26755 41599
rect 28074 41596 28080 41608
rect 26743 41568 28080 41596
rect 26743 41565 26755 41568
rect 26697 41559 26755 41565
rect 28074 41556 28080 41568
rect 28132 41556 28138 41608
rect 28629 41599 28687 41605
rect 28629 41565 28641 41599
rect 28675 41565 28687 41599
rect 28629 41559 28687 41565
rect 23382 41488 23388 41540
rect 23440 41528 23446 41540
rect 24826 41531 24884 41537
rect 24826 41528 24838 41531
rect 23440 41500 24838 41528
rect 23440 41488 23446 41500
rect 24826 41497 24838 41500
rect 24872 41497 24884 41531
rect 24826 41491 24884 41497
rect 26964 41531 27022 41537
rect 26964 41497 26976 41531
rect 27010 41528 27022 41531
rect 27338 41528 27344 41540
rect 27010 41500 27344 41528
rect 27010 41497 27022 41500
rect 26964 41491 27022 41497
rect 27338 41488 27344 41500
rect 27396 41488 27402 41540
rect 28644 41528 28672 41559
rect 28718 41556 28724 41608
rect 28776 41596 28782 41608
rect 28776 41568 28821 41596
rect 28776 41556 28782 41568
rect 30558 41556 30564 41608
rect 30616 41596 30622 41608
rect 30745 41599 30803 41605
rect 30745 41596 30757 41599
rect 30616 41568 30757 41596
rect 30616 41556 30622 41568
rect 30745 41565 30757 41568
rect 30791 41565 30803 41599
rect 31573 41599 31631 41605
rect 30745 41559 30803 41565
rect 30852 41568 31248 41596
rect 29914 41528 29920 41540
rect 28644 41500 29920 41528
rect 29914 41488 29920 41500
rect 29972 41488 29978 41540
rect 30650 41488 30656 41540
rect 30708 41528 30714 41540
rect 30852 41537 30880 41568
rect 30837 41531 30895 41537
rect 30837 41528 30849 41531
rect 30708 41500 30849 41528
rect 30708 41488 30714 41500
rect 30837 41497 30849 41500
rect 30883 41497 30895 41531
rect 30837 41491 30895 41497
rect 31018 41488 31024 41540
rect 31076 41528 31082 41540
rect 31113 41531 31171 41537
rect 31113 41528 31125 41531
rect 31076 41500 31125 41528
rect 31076 41488 31082 41500
rect 31113 41497 31125 41500
rect 31159 41497 31171 41531
rect 31113 41491 31171 41497
rect 30926 41420 30932 41472
rect 30984 41460 30990 41472
rect 31220 41460 31248 41568
rect 31573 41565 31585 41599
rect 31619 41596 31631 41599
rect 32122 41596 32128 41608
rect 31619 41568 32128 41596
rect 31619 41565 31631 41568
rect 31573 41559 31631 41565
rect 32122 41556 32128 41568
rect 32180 41556 32186 41608
rect 34790 41556 34796 41608
rect 34848 41596 34854 41608
rect 34885 41599 34943 41605
rect 34885 41596 34897 41599
rect 34848 41568 34897 41596
rect 34848 41556 34854 41568
rect 34885 41565 34897 41568
rect 34931 41565 34943 41599
rect 34885 41559 34943 41565
rect 35069 41599 35127 41605
rect 35069 41565 35081 41599
rect 35115 41596 35127 41599
rect 35866 41596 35894 41760
rect 38194 41664 38200 41676
rect 38155 41636 38200 41664
rect 38194 41624 38200 41636
rect 38252 41624 38258 41676
rect 43162 41664 43168 41676
rect 42720 41636 43168 41664
rect 35115 41568 35894 41596
rect 36357 41599 36415 41605
rect 35115 41565 35127 41568
rect 35069 41559 35127 41565
rect 36357 41565 36369 41599
rect 36403 41596 36415 41599
rect 37458 41596 37464 41608
rect 36403 41568 37464 41596
rect 36403 41565 36415 41568
rect 36357 41559 36415 41565
rect 31840 41531 31898 41537
rect 31840 41497 31852 41531
rect 31886 41528 31898 41531
rect 32306 41528 32312 41540
rect 31886 41500 32312 41528
rect 31886 41497 31898 41500
rect 31840 41491 31898 41497
rect 32306 41488 32312 41500
rect 32364 41488 32370 41540
rect 34054 41488 34060 41540
rect 34112 41528 34118 41540
rect 35084 41528 35112 41559
rect 37458 41556 37464 41568
rect 37516 41556 37522 41608
rect 37642 41556 37648 41608
rect 37700 41596 37706 41608
rect 42720 41605 42748 41636
rect 43162 41624 43168 41636
rect 43220 41624 43226 41676
rect 46474 41664 46480 41676
rect 46435 41636 46480 41664
rect 46474 41624 46480 41636
rect 46532 41624 46538 41676
rect 46661 41667 46719 41673
rect 46661 41633 46673 41667
rect 46707 41664 46719 41667
rect 47854 41664 47860 41676
rect 46707 41636 47860 41664
rect 46707 41633 46719 41636
rect 46661 41627 46719 41633
rect 47854 41624 47860 41636
rect 47912 41624 47918 41676
rect 48222 41664 48228 41676
rect 48183 41636 48228 41664
rect 48222 41624 48228 41636
rect 48280 41624 48286 41676
rect 38381 41599 38439 41605
rect 38381 41596 38393 41599
rect 37700 41568 38393 41596
rect 37700 41556 37706 41568
rect 38381 41565 38393 41568
rect 38427 41565 38439 41599
rect 38381 41559 38439 41565
rect 42705 41599 42763 41605
rect 42705 41565 42717 41599
rect 42751 41565 42763 41599
rect 42705 41559 42763 41565
rect 42886 41556 42892 41608
rect 42944 41596 42950 41608
rect 43073 41599 43131 41605
rect 42944 41568 43037 41596
rect 42944 41556 42950 41568
rect 34112 41500 35112 41528
rect 36624 41531 36682 41537
rect 34112 41488 34118 41500
rect 36624 41497 36636 41531
rect 36670 41528 36682 41531
rect 36722 41528 36728 41540
rect 36670 41500 36728 41528
rect 36670 41497 36682 41500
rect 36624 41491 36682 41497
rect 36722 41488 36728 41500
rect 36780 41488 36786 41540
rect 42996 41528 43024 41568
rect 43073 41565 43085 41599
rect 43119 41596 43131 41599
rect 43717 41599 43775 41605
rect 43717 41596 43729 41599
rect 43119 41568 43729 41596
rect 43119 41565 43131 41568
rect 43073 41559 43131 41565
rect 43717 41565 43729 41568
rect 43763 41565 43775 41599
rect 43717 41559 43775 41565
rect 45373 41599 45431 41605
rect 45373 41565 45385 41599
rect 45419 41596 45431 41599
rect 45554 41596 45560 41608
rect 45419 41568 45560 41596
rect 45419 41565 45431 41568
rect 45373 41559 45431 41565
rect 45554 41556 45560 41568
rect 45612 41556 45618 41608
rect 44082 41528 44088 41540
rect 42996 41500 44088 41528
rect 44082 41488 44088 41500
rect 44140 41488 44146 41540
rect 32953 41463 33011 41469
rect 32953 41460 32965 41463
rect 30984 41432 31029 41460
rect 31220 41432 32965 41460
rect 30984 41420 30990 41432
rect 32953 41429 32965 41432
rect 32999 41429 33011 41463
rect 37734 41460 37740 41472
rect 37647 41432 37740 41460
rect 32953 41423 33011 41429
rect 37734 41420 37740 41432
rect 37792 41460 37798 41472
rect 38194 41460 38200 41472
rect 37792 41432 38200 41460
rect 37792 41420 37798 41432
rect 38194 41420 38200 41432
rect 38252 41420 38258 41472
rect 45186 41460 45192 41472
rect 45147 41432 45192 41460
rect 45186 41420 45192 41432
rect 45244 41420 45250 41472
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 32490 41216 32496 41268
rect 32548 41256 32554 41268
rect 32677 41259 32735 41265
rect 32677 41256 32689 41259
rect 32548 41228 32689 41256
rect 32548 41216 32554 41228
rect 32677 41225 32689 41228
rect 32723 41225 32735 41259
rect 32677 41219 32735 41225
rect 33134 41216 33140 41268
rect 33192 41256 33198 41268
rect 34054 41256 34060 41268
rect 33192 41228 34060 41256
rect 33192 41216 33198 41228
rect 34054 41216 34060 41228
rect 34112 41216 34118 41268
rect 35618 41216 35624 41268
rect 35676 41256 35682 41268
rect 35676 41228 47808 41256
rect 35676 41216 35682 41228
rect 30561 41191 30619 41197
rect 30561 41157 30573 41191
rect 30607 41188 30619 41191
rect 30926 41188 30932 41200
rect 30607 41160 30932 41188
rect 30607 41157 30619 41160
rect 30561 41151 30619 41157
rect 30926 41148 30932 41160
rect 30984 41188 30990 41200
rect 30984 41160 31754 41188
rect 30984 41148 30990 41160
rect 2038 41120 2044 41132
rect 1999 41092 2044 41120
rect 2038 41080 2044 41092
rect 2096 41080 2102 41132
rect 24213 41123 24271 41129
rect 24213 41089 24225 41123
rect 24259 41120 24271 41123
rect 24302 41120 24308 41132
rect 24259 41092 24308 41120
rect 24259 41089 24271 41092
rect 24213 41083 24271 41089
rect 24302 41080 24308 41092
rect 24360 41080 24366 41132
rect 24486 41129 24492 41132
rect 24480 41083 24492 41129
rect 24544 41120 24550 41132
rect 30837 41123 30895 41129
rect 24544 41092 24580 41120
rect 24486 41080 24492 41083
rect 24544 41080 24550 41092
rect 30837 41089 30849 41123
rect 30883 41120 30895 41123
rect 31110 41120 31116 41132
rect 30883 41092 31116 41120
rect 30883 41089 30895 41092
rect 30837 41083 30895 41089
rect 31110 41080 31116 41092
rect 31168 41080 31174 41132
rect 31726 41120 31754 41160
rect 32398 41120 32404 41132
rect 31726 41092 32404 41120
rect 32398 41080 32404 41092
rect 32456 41080 32462 41132
rect 32493 41123 32551 41129
rect 32493 41089 32505 41123
rect 32539 41120 32551 41123
rect 33152 41120 33180 41216
rect 37366 41148 37372 41200
rect 37424 41188 37430 41200
rect 37424 41160 38240 41188
rect 37424 41148 37430 41160
rect 33962 41120 33968 41132
rect 32539 41092 33180 41120
rect 33923 41092 33968 41120
rect 32539 41089 32551 41092
rect 32493 41083 32551 41089
rect 33962 41080 33968 41092
rect 34020 41080 34026 41132
rect 36449 41123 36507 41129
rect 36449 41089 36461 41123
rect 36495 41120 36507 41123
rect 36725 41123 36783 41129
rect 36495 41092 36676 41120
rect 36495 41089 36507 41092
rect 36449 41083 36507 41089
rect 2225 41055 2283 41061
rect 2225 41021 2237 41055
rect 2271 41052 2283 41055
rect 2406 41052 2412 41064
rect 2271 41024 2412 41052
rect 2271 41021 2283 41024
rect 2225 41015 2283 41021
rect 2406 41012 2412 41024
rect 2464 41012 2470 41064
rect 2774 41052 2780 41064
rect 2735 41024 2780 41052
rect 2774 41012 2780 41024
rect 2832 41012 2838 41064
rect 30650 41052 30656 41064
rect 30611 41024 30656 41052
rect 30650 41012 30656 41024
rect 30708 41012 30714 41064
rect 36538 41052 36544 41064
rect 36499 41024 36544 41052
rect 36538 41012 36544 41024
rect 36596 41012 36602 41064
rect 36648 41052 36676 41092
rect 36725 41089 36737 41123
rect 36771 41120 36783 41123
rect 37274 41120 37280 41132
rect 36771 41092 37280 41120
rect 36771 41089 36783 41092
rect 36725 41083 36783 41089
rect 37274 41080 37280 41092
rect 37332 41120 37338 41132
rect 37734 41120 37740 41132
rect 37332 41092 37740 41120
rect 37332 41080 37338 41092
rect 37734 41080 37740 41092
rect 37792 41080 37798 41132
rect 38212 41120 38240 41160
rect 38286 41148 38292 41200
rect 38344 41188 38350 41200
rect 38442 41191 38500 41197
rect 38442 41188 38454 41191
rect 38344 41160 38454 41188
rect 38344 41148 38350 41160
rect 38442 41157 38454 41160
rect 38488 41157 38500 41191
rect 42886 41188 42892 41200
rect 38442 41151 38500 41157
rect 41892 41160 42892 41188
rect 40218 41120 40224 41132
rect 38212 41092 39620 41120
rect 40179 41092 40224 41120
rect 37366 41052 37372 41064
rect 36648 41024 37372 41052
rect 37366 41012 37372 41024
rect 37424 41012 37430 41064
rect 37458 41012 37464 41064
rect 37516 41052 37522 41064
rect 38197 41055 38255 41061
rect 38197 41052 38209 41055
rect 37516 41024 38209 41052
rect 37516 41012 37522 41024
rect 38197 41021 38209 41024
rect 38243 41021 38255 41055
rect 38197 41015 38255 41021
rect 37182 40984 37188 40996
rect 36556 40956 37188 40984
rect 25590 40916 25596 40928
rect 25551 40888 25596 40916
rect 25590 40876 25596 40888
rect 25648 40876 25654 40928
rect 30558 40916 30564 40928
rect 30519 40888 30564 40916
rect 30558 40876 30564 40888
rect 30616 40876 30622 40928
rect 30834 40876 30840 40928
rect 30892 40916 30898 40928
rect 31021 40919 31079 40925
rect 31021 40916 31033 40919
rect 30892 40888 31033 40916
rect 30892 40876 30898 40888
rect 31021 40885 31033 40888
rect 31067 40885 31079 40919
rect 33778 40916 33784 40928
rect 33739 40888 33784 40916
rect 31021 40879 31079 40885
rect 33778 40876 33784 40888
rect 33836 40876 33842 40928
rect 36556 40925 36584 40956
rect 37182 40944 37188 40956
rect 37240 40944 37246 40996
rect 36541 40919 36599 40925
rect 36541 40885 36553 40919
rect 36587 40885 36599 40919
rect 36541 40879 36599 40885
rect 36630 40876 36636 40928
rect 36688 40916 36694 40928
rect 36909 40919 36967 40925
rect 36909 40916 36921 40919
rect 36688 40888 36921 40916
rect 36688 40876 36694 40888
rect 36909 40885 36921 40888
rect 36955 40885 36967 40919
rect 38212 40916 38240 41015
rect 39592 40996 39620 41092
rect 40218 41080 40224 41092
rect 40276 41080 40282 41132
rect 41233 41123 41291 41129
rect 41233 41089 41245 41123
rect 41279 41120 41291 41123
rect 41782 41120 41788 41132
rect 41279 41092 41788 41120
rect 41279 41089 41291 41092
rect 41233 41083 41291 41089
rect 41782 41080 41788 41092
rect 41840 41080 41846 41132
rect 41892 41129 41920 41160
rect 42886 41148 42892 41160
rect 42944 41148 42950 41200
rect 44904 41191 44962 41197
rect 44904 41157 44916 41191
rect 44950 41188 44962 41191
rect 45186 41188 45192 41200
rect 44950 41160 45192 41188
rect 44950 41157 44962 41160
rect 44904 41151 44962 41157
rect 45186 41148 45192 41160
rect 45244 41148 45250 41200
rect 41877 41123 41935 41129
rect 41877 41089 41889 41123
rect 41923 41089 41935 41123
rect 42797 41123 42855 41129
rect 42797 41120 42809 41123
rect 41877 41083 41935 41089
rect 42720 41092 42809 41120
rect 41693 41055 41751 41061
rect 41693 41021 41705 41055
rect 41739 41052 41751 41055
rect 42242 41052 42248 41064
rect 41739 41024 42248 41052
rect 41739 41021 41751 41024
rect 41693 41015 41751 41021
rect 42242 41012 42248 41024
rect 42300 41052 42306 41064
rect 42720 41052 42748 41092
rect 42797 41089 42809 41092
rect 42843 41089 42855 41123
rect 43070 41120 43076 41132
rect 42983 41092 43076 41120
rect 42797 41083 42855 41089
rect 43070 41080 43076 41092
rect 43128 41120 43134 41132
rect 43990 41120 43996 41132
rect 43128 41092 43996 41120
rect 43128 41080 43134 41092
rect 43990 41080 43996 41092
rect 44048 41080 44054 41132
rect 44637 41123 44695 41129
rect 44637 41089 44649 41123
rect 44683 41120 44695 41123
rect 44726 41120 44732 41132
rect 44683 41092 44732 41120
rect 44683 41089 44695 41092
rect 44637 41083 44695 41089
rect 44726 41080 44732 41092
rect 44784 41080 44790 41132
rect 47780 41129 47808 41228
rect 47765 41123 47823 41129
rect 47765 41089 47777 41123
rect 47811 41089 47823 41123
rect 47765 41083 47823 41089
rect 42886 41052 42892 41064
rect 42300 41024 42748 41052
rect 42847 41024 42892 41052
rect 42300 41012 42306 41024
rect 42886 41012 42892 41024
rect 42944 41012 42950 41064
rect 39574 40984 39580 40996
rect 39487 40956 39580 40984
rect 39574 40944 39580 40956
rect 39632 40944 39638 40996
rect 43162 40984 43168 40996
rect 43075 40956 43168 40984
rect 38562 40916 38568 40928
rect 38212 40888 38568 40916
rect 36909 40879 36967 40885
rect 38562 40876 38568 40888
rect 38620 40876 38626 40928
rect 39666 40876 39672 40928
rect 39724 40916 39730 40928
rect 40037 40919 40095 40925
rect 40037 40916 40049 40919
rect 39724 40888 40049 40916
rect 39724 40876 39730 40888
rect 40037 40885 40049 40888
rect 40083 40885 40095 40919
rect 40037 40879 40095 40885
rect 41049 40919 41107 40925
rect 41049 40885 41061 40919
rect 41095 40916 41107 40919
rect 41138 40916 41144 40928
rect 41095 40888 41144 40916
rect 41095 40885 41107 40888
rect 41049 40879 41107 40885
rect 41138 40876 41144 40888
rect 41196 40876 41202 40928
rect 42061 40919 42119 40925
rect 42061 40885 42073 40919
rect 42107 40916 42119 40919
rect 42518 40916 42524 40928
rect 42107 40888 42524 40916
rect 42107 40885 42119 40888
rect 42061 40879 42119 40885
rect 42518 40876 42524 40888
rect 42576 40876 42582 40928
rect 43088 40925 43116 40956
rect 43162 40944 43168 40956
rect 43220 40984 43226 40996
rect 43220 40956 43484 40984
rect 43220 40944 43226 40956
rect 43073 40919 43131 40925
rect 43073 40885 43085 40919
rect 43119 40885 43131 40919
rect 43254 40916 43260 40928
rect 43215 40888 43260 40916
rect 43073 40879 43131 40885
rect 43254 40876 43260 40888
rect 43312 40876 43318 40928
rect 43456 40916 43484 40956
rect 46017 40919 46075 40925
rect 46017 40916 46029 40919
rect 43456 40888 46029 40916
rect 46017 40885 46029 40888
rect 46063 40885 46075 40919
rect 46017 40879 46075 40885
rect 46474 40876 46480 40928
rect 46532 40916 46538 40928
rect 47213 40919 47271 40925
rect 47213 40916 47225 40919
rect 46532 40888 47225 40916
rect 46532 40876 46538 40888
rect 47213 40885 47225 40888
rect 47259 40885 47271 40919
rect 47854 40916 47860 40928
rect 47815 40888 47860 40916
rect 47213 40879 47271 40885
rect 47854 40876 47860 40888
rect 47912 40876 47918 40928
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 2406 40712 2412 40724
rect 2367 40684 2412 40712
rect 2406 40672 2412 40684
rect 2464 40672 2470 40724
rect 23845 40715 23903 40721
rect 23845 40681 23857 40715
rect 23891 40712 23903 40715
rect 24486 40712 24492 40724
rect 23891 40684 24492 40712
rect 23891 40681 23903 40684
rect 23845 40675 23903 40681
rect 24486 40672 24492 40684
rect 24544 40672 24550 40724
rect 28258 40672 28264 40724
rect 28316 40712 28322 40724
rect 28534 40712 28540 40724
rect 28316 40684 28540 40712
rect 28316 40672 28322 40684
rect 28534 40672 28540 40684
rect 28592 40672 28598 40724
rect 29914 40712 29920 40724
rect 29875 40684 29920 40712
rect 29914 40672 29920 40684
rect 29972 40672 29978 40724
rect 34333 40715 34391 40721
rect 34333 40681 34345 40715
rect 34379 40712 34391 40715
rect 34790 40712 34796 40724
rect 34379 40684 34796 40712
rect 34379 40681 34391 40684
rect 34333 40675 34391 40681
rect 34790 40672 34796 40684
rect 34848 40712 34854 40724
rect 35713 40715 35771 40721
rect 35713 40712 35725 40715
rect 34848 40684 35725 40712
rect 34848 40672 34854 40684
rect 35713 40681 35725 40684
rect 35759 40712 35771 40715
rect 35802 40712 35808 40724
rect 35759 40684 35808 40712
rect 35759 40681 35771 40684
rect 35713 40675 35771 40681
rect 35802 40672 35808 40684
rect 35860 40672 35866 40724
rect 42242 40712 42248 40724
rect 42203 40684 42248 40712
rect 42242 40672 42248 40684
rect 42300 40672 42306 40724
rect 45554 40712 45560 40724
rect 45515 40684 45560 40712
rect 45554 40672 45560 40684
rect 45612 40672 45618 40724
rect 28626 40604 28632 40656
rect 28684 40604 28690 40656
rect 36909 40647 36967 40653
rect 36909 40613 36921 40647
rect 36955 40644 36967 40647
rect 37274 40644 37280 40656
rect 36955 40616 37280 40644
rect 36955 40613 36967 40616
rect 36909 40607 36967 40613
rect 37274 40604 37280 40616
rect 37332 40604 37338 40656
rect 24949 40579 25007 40585
rect 24949 40576 24961 40579
rect 24044 40548 24961 40576
rect 2222 40468 2228 40520
rect 2280 40508 2286 40520
rect 2317 40511 2375 40517
rect 2317 40508 2329 40511
rect 2280 40480 2329 40508
rect 2280 40468 2286 40480
rect 2317 40477 2329 40480
rect 2363 40508 2375 40511
rect 4706 40508 4712 40520
rect 2363 40480 4712 40508
rect 2363 40477 2375 40480
rect 2317 40471 2375 40477
rect 4706 40468 4712 40480
rect 4764 40468 4770 40520
rect 24044 40517 24072 40548
rect 24949 40545 24961 40548
rect 24995 40545 25007 40579
rect 28644 40576 28672 40604
rect 24949 40539 25007 40545
rect 28552 40548 28672 40576
rect 24029 40511 24087 40517
rect 24029 40477 24041 40511
rect 24075 40477 24087 40511
rect 24029 40471 24087 40477
rect 24673 40511 24731 40517
rect 24673 40477 24685 40511
rect 24719 40477 24731 40511
rect 24673 40471 24731 40477
rect 24688 40440 24716 40471
rect 24762 40468 24768 40520
rect 24820 40508 24826 40520
rect 28552 40517 28580 40548
rect 32122 40536 32128 40588
rect 32180 40576 32186 40588
rect 32950 40576 32956 40588
rect 32180 40548 32956 40576
rect 32180 40536 32186 40548
rect 32950 40536 32956 40548
rect 33008 40536 33014 40588
rect 38562 40536 38568 40588
rect 38620 40576 38626 40588
rect 40865 40579 40923 40585
rect 40865 40576 40877 40579
rect 38620 40548 40877 40576
rect 38620 40536 38626 40548
rect 40865 40545 40877 40548
rect 40911 40545 40923 40579
rect 40865 40539 40923 40545
rect 44082 40536 44088 40588
rect 44140 40576 44146 40588
rect 46474 40576 46480 40588
rect 44140 40548 45416 40576
rect 46435 40548 46480 40576
rect 44140 40536 44146 40548
rect 28537 40511 28595 40517
rect 24820 40480 24865 40508
rect 24820 40468 24826 40480
rect 28537 40477 28549 40511
rect 28583 40477 28595 40511
rect 28537 40471 28595 40477
rect 28721 40511 28779 40517
rect 28721 40477 28733 40511
rect 28767 40508 28779 40511
rect 33220 40511 33278 40517
rect 28767 40480 29776 40508
rect 28767 40477 28779 40480
rect 28721 40471 28779 40477
rect 29748 40452 29776 40480
rect 33220 40477 33232 40511
rect 33266 40508 33278 40511
rect 33778 40508 33784 40520
rect 33266 40480 33784 40508
rect 33266 40477 33278 40480
rect 33220 40471 33278 40477
rect 33778 40468 33784 40480
rect 33836 40468 33842 40520
rect 37461 40511 37519 40517
rect 37461 40508 37473 40511
rect 36639 40480 37473 40508
rect 25038 40440 25044 40452
rect 24688 40412 25044 40440
rect 25038 40400 25044 40412
rect 25096 40400 25102 40452
rect 29730 40440 29736 40452
rect 29643 40412 29736 40440
rect 29730 40400 29736 40412
rect 29788 40400 29794 40452
rect 29949 40443 30007 40449
rect 29949 40409 29961 40443
rect 29995 40440 30007 40443
rect 31018 40440 31024 40452
rect 29995 40412 31024 40440
rect 29995 40409 30007 40412
rect 29949 40403 30007 40409
rect 31018 40400 31024 40412
rect 31076 40400 31082 40452
rect 34514 40400 34520 40452
rect 34572 40440 34578 40452
rect 35529 40443 35587 40449
rect 35529 40440 35541 40443
rect 34572 40412 35541 40440
rect 34572 40400 34578 40412
rect 35529 40409 35541 40412
rect 35575 40409 35587 40443
rect 35529 40403 35587 40409
rect 35745 40443 35803 40449
rect 35745 40409 35757 40443
rect 35791 40440 35803 40443
rect 36639 40440 36667 40480
rect 37461 40477 37473 40480
rect 37507 40477 37519 40511
rect 37461 40471 37519 40477
rect 39393 40511 39451 40517
rect 39393 40477 39405 40511
rect 39439 40477 39451 40511
rect 39393 40471 39451 40477
rect 37090 40440 37096 40452
rect 35791 40412 36667 40440
rect 37051 40412 37096 40440
rect 35791 40409 35803 40412
rect 35745 40403 35803 40409
rect 37090 40400 37096 40412
rect 37148 40400 37154 40452
rect 37277 40443 37335 40449
rect 37277 40409 37289 40443
rect 37323 40440 37335 40443
rect 37366 40440 37372 40452
rect 37323 40412 37372 40440
rect 37323 40409 37335 40412
rect 37277 40403 37335 40409
rect 37366 40400 37372 40412
rect 37424 40400 37430 40452
rect 39408 40440 39436 40471
rect 39574 40468 39580 40520
rect 39632 40508 39638 40520
rect 40037 40511 40095 40517
rect 40037 40508 40049 40511
rect 39632 40480 40049 40508
rect 39632 40468 39638 40480
rect 40037 40477 40049 40480
rect 40083 40477 40095 40511
rect 40218 40508 40224 40520
rect 40179 40480 40224 40508
rect 40037 40471 40095 40477
rect 40218 40468 40224 40480
rect 40276 40508 40282 40520
rect 41138 40517 41144 40520
rect 41132 40508 41144 40517
rect 40276 40480 40540 40508
rect 41099 40480 41144 40508
rect 40276 40468 40282 40480
rect 40405 40443 40463 40449
rect 40405 40440 40417 40443
rect 39408 40412 40417 40440
rect 40405 40409 40417 40412
rect 40451 40409 40463 40443
rect 40512 40440 40540 40480
rect 41132 40471 41144 40480
rect 41138 40468 41144 40471
rect 41196 40468 41202 40520
rect 42610 40468 42616 40520
rect 42668 40508 42674 40520
rect 42705 40511 42763 40517
rect 42705 40508 42717 40511
rect 42668 40480 42717 40508
rect 42668 40468 42674 40480
rect 42705 40477 42717 40480
rect 42751 40508 42763 40511
rect 44726 40508 44732 40520
rect 42751 40480 44732 40508
rect 42751 40477 42763 40480
rect 42705 40471 42763 40477
rect 44726 40468 44732 40480
rect 44784 40468 44790 40520
rect 45278 40508 45284 40520
rect 45239 40480 45284 40508
rect 45278 40468 45284 40480
rect 45336 40468 45342 40520
rect 45388 40517 45416 40548
rect 46474 40536 46480 40548
rect 46532 40536 46538 40588
rect 46661 40579 46719 40585
rect 46661 40545 46673 40579
rect 46707 40576 46719 40579
rect 47854 40576 47860 40588
rect 46707 40548 47860 40576
rect 46707 40545 46719 40548
rect 46661 40539 46719 40545
rect 47854 40536 47860 40548
rect 47912 40536 47918 40588
rect 48222 40576 48228 40588
rect 48183 40548 48228 40576
rect 48222 40536 48228 40548
rect 48280 40536 48286 40588
rect 45373 40511 45431 40517
rect 45373 40477 45385 40511
rect 45419 40477 45431 40511
rect 45373 40471 45431 40477
rect 41598 40440 41604 40452
rect 40512 40412 41604 40440
rect 40405 40403 40463 40409
rect 41598 40400 41604 40412
rect 41656 40440 41662 40452
rect 42794 40440 42800 40452
rect 41656 40412 42800 40440
rect 41656 40400 41662 40412
rect 42794 40400 42800 40412
rect 42852 40400 42858 40452
rect 42978 40449 42984 40452
rect 42972 40403 42984 40449
rect 43036 40440 43042 40452
rect 43036 40412 43072 40440
rect 42978 40400 42984 40403
rect 43036 40400 43042 40412
rect 28905 40375 28963 40381
rect 28905 40341 28917 40375
rect 28951 40372 28963 40375
rect 29822 40372 29828 40384
rect 28951 40344 29828 40372
rect 28951 40341 28963 40344
rect 28905 40335 28963 40341
rect 29822 40332 29828 40344
rect 29880 40332 29886 40384
rect 30098 40372 30104 40384
rect 30059 40344 30104 40372
rect 30098 40332 30104 40344
rect 30156 40332 30162 40384
rect 35342 40332 35348 40384
rect 35400 40372 35406 40384
rect 35897 40375 35955 40381
rect 35897 40372 35909 40375
rect 35400 40344 35909 40372
rect 35400 40332 35406 40344
rect 35897 40341 35909 40344
rect 35943 40341 35955 40375
rect 35897 40335 35955 40341
rect 36538 40332 36544 40384
rect 36596 40372 36602 40384
rect 37182 40372 37188 40384
rect 36596 40344 37188 40372
rect 36596 40332 36602 40344
rect 37182 40332 37188 40344
rect 37240 40332 37246 40384
rect 39206 40372 39212 40384
rect 39167 40344 39212 40372
rect 39206 40332 39212 40344
rect 39264 40332 39270 40384
rect 42886 40332 42892 40384
rect 42944 40372 42950 40384
rect 44085 40375 44143 40381
rect 44085 40372 44097 40375
rect 42944 40344 44097 40372
rect 42944 40332 42950 40344
rect 44085 40341 44097 40344
rect 44131 40341 44143 40375
rect 44085 40335 44143 40341
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 25038 40168 25044 40180
rect 24999 40140 25044 40168
rect 25038 40128 25044 40140
rect 25096 40128 25102 40180
rect 27985 40171 28043 40177
rect 27985 40137 27997 40171
rect 28031 40137 28043 40171
rect 27985 40131 28043 40137
rect 28000 40100 28028 40131
rect 29914 40128 29920 40180
rect 29972 40168 29978 40180
rect 30009 40171 30067 40177
rect 30009 40168 30021 40171
rect 29972 40140 30021 40168
rect 29972 40128 29978 40140
rect 30009 40137 30021 40140
rect 30055 40137 30067 40171
rect 34514 40168 34520 40180
rect 34475 40140 34520 40168
rect 30009 40131 30067 40137
rect 28874 40103 28932 40109
rect 28874 40100 28886 40103
rect 28000 40072 28886 40100
rect 28874 40069 28886 40072
rect 28920 40069 28932 40103
rect 30024 40100 30052 40131
rect 34514 40128 34520 40140
rect 34572 40128 34578 40180
rect 35802 40128 35808 40180
rect 35860 40168 35866 40180
rect 35860 40140 36492 40168
rect 35860 40128 35866 40140
rect 30024 40072 30696 40100
rect 28874 40063 28932 40069
rect 23934 40041 23940 40044
rect 23928 39995 23940 40041
rect 23992 40032 23998 40044
rect 25590 40032 25596 40044
rect 23992 40004 24028 40032
rect 25551 40004 25596 40032
rect 23934 39992 23940 39995
rect 23992 39992 23998 40004
rect 25590 39992 25596 40004
rect 25648 39992 25654 40044
rect 25777 40035 25835 40041
rect 25777 40001 25789 40035
rect 25823 40032 25835 40035
rect 28169 40035 28227 40041
rect 25823 40004 27292 40032
rect 25823 40001 25835 40004
rect 25777 39995 25835 40001
rect 23661 39967 23719 39973
rect 23661 39933 23673 39967
rect 23707 39933 23719 39967
rect 23661 39927 23719 39933
rect 23676 39828 23704 39927
rect 24762 39924 24768 39976
rect 24820 39964 24826 39976
rect 25792 39964 25820 39995
rect 24820 39936 25820 39964
rect 24820 39924 24826 39936
rect 24302 39828 24308 39840
rect 23676 39800 24308 39828
rect 24302 39788 24308 39800
rect 24360 39828 24366 39840
rect 24578 39828 24584 39840
rect 24360 39800 24584 39828
rect 24360 39788 24366 39800
rect 24578 39788 24584 39800
rect 24636 39788 24642 39840
rect 25961 39831 26019 39837
rect 25961 39797 25973 39831
rect 26007 39828 26019 39831
rect 26602 39828 26608 39840
rect 26007 39800 26608 39828
rect 26007 39797 26019 39800
rect 25961 39791 26019 39797
rect 26602 39788 26608 39800
rect 26660 39788 26666 39840
rect 27264 39828 27292 40004
rect 28169 40001 28181 40035
rect 28215 40032 28227 40035
rect 30006 40032 30012 40044
rect 28215 40004 30012 40032
rect 28215 40001 28227 40004
rect 28169 39995 28227 40001
rect 30006 39992 30012 40004
rect 30064 39992 30070 40044
rect 30668 40041 30696 40072
rect 33888 40072 35296 40100
rect 30653 40035 30711 40041
rect 30653 40001 30665 40035
rect 30699 40001 30711 40035
rect 30834 40032 30840 40044
rect 30795 40004 30840 40032
rect 30653 39995 30711 40001
rect 30834 39992 30840 40004
rect 30892 39992 30898 40044
rect 30926 39992 30932 40044
rect 30984 40032 30990 40044
rect 30984 40004 31029 40032
rect 30984 39992 30990 40004
rect 32950 39992 32956 40044
rect 33008 40032 33014 40044
rect 33137 40035 33195 40041
rect 33137 40032 33149 40035
rect 33008 40004 33149 40032
rect 33008 39992 33014 40004
rect 33137 40001 33149 40004
rect 33183 40001 33195 40035
rect 33137 39995 33195 40001
rect 33226 39992 33232 40044
rect 33284 40032 33290 40044
rect 33404 40035 33462 40041
rect 33404 40032 33416 40035
rect 33284 40004 33416 40032
rect 33284 39992 33290 40004
rect 33404 40001 33416 40004
rect 33450 40032 33462 40035
rect 33888 40032 33916 40072
rect 33450 40004 33916 40032
rect 33450 40001 33462 40004
rect 33404 39995 33462 40001
rect 28074 39924 28080 39976
rect 28132 39964 28138 39976
rect 28629 39967 28687 39973
rect 28629 39964 28641 39967
rect 28132 39936 28641 39964
rect 28132 39924 28138 39936
rect 28629 39933 28641 39936
rect 28675 39933 28687 39967
rect 28629 39927 28687 39933
rect 29822 39924 29828 39976
rect 29880 39964 29886 39976
rect 30745 39967 30803 39973
rect 30745 39964 30757 39967
rect 29880 39936 30757 39964
rect 29880 39924 29886 39936
rect 30745 39933 30757 39936
rect 30791 39933 30803 39967
rect 35268 39964 35296 40072
rect 35342 40060 35348 40112
rect 35400 40060 35406 40112
rect 35526 40100 35532 40112
rect 35487 40072 35532 40100
rect 35526 40060 35532 40072
rect 35584 40060 35590 40112
rect 35667 40103 35725 40109
rect 35667 40069 35679 40103
rect 35713 40100 35725 40103
rect 36265 40103 36323 40109
rect 36265 40100 36277 40103
rect 35713 40072 36277 40100
rect 35713 40069 35725 40072
rect 35667 40063 35725 40069
rect 36265 40069 36277 40072
rect 36311 40069 36323 40103
rect 36265 40063 36323 40069
rect 35346 40057 35404 40060
rect 35346 40023 35358 40057
rect 35392 40023 35404 40057
rect 36464 40041 36492 40140
rect 37182 40128 37188 40180
rect 37240 40168 37246 40180
rect 40037 40171 40095 40177
rect 40037 40168 40049 40171
rect 37240 40140 40049 40168
rect 37240 40128 37246 40140
rect 40037 40137 40049 40140
rect 40083 40137 40095 40171
rect 42886 40168 42892 40180
rect 42847 40140 42892 40168
rect 40037 40131 40095 40137
rect 42886 40128 42892 40140
rect 42944 40128 42950 40180
rect 45278 40128 45284 40180
rect 45336 40168 45342 40180
rect 46109 40171 46167 40177
rect 46109 40168 46121 40171
rect 45336 40140 46121 40168
rect 45336 40128 45342 40140
rect 46109 40137 46121 40140
rect 46155 40137 46167 40171
rect 46109 40131 46167 40137
rect 38924 40103 38982 40109
rect 38924 40069 38936 40103
rect 38970 40100 38982 40103
rect 39206 40100 39212 40112
rect 38970 40072 39212 40100
rect 38970 40069 38982 40072
rect 38924 40063 38982 40069
rect 39206 40060 39212 40072
rect 39264 40060 39270 40112
rect 42242 40060 42248 40112
rect 42300 40100 42306 40112
rect 42981 40103 43039 40109
rect 42981 40100 42993 40103
rect 42300 40072 42993 40100
rect 42300 40060 42306 40072
rect 42981 40069 42993 40072
rect 43027 40069 43039 40103
rect 43162 40100 43168 40112
rect 42981 40063 43039 40069
rect 43088 40072 43168 40100
rect 35346 40017 35404 40023
rect 35437 40035 35495 40041
rect 35437 40001 35449 40035
rect 35483 40001 35495 40035
rect 35437 39995 35495 40001
rect 36449 40035 36507 40041
rect 36449 40001 36461 40035
rect 36495 40001 36507 40035
rect 36630 40032 36636 40044
rect 36591 40004 36636 40032
rect 36449 39995 36507 40001
rect 35452 39964 35480 39995
rect 36630 39992 36636 40004
rect 36688 39992 36694 40044
rect 36722 39992 36728 40044
rect 36780 40032 36786 40044
rect 41598 40032 41604 40044
rect 36780 40004 36825 40032
rect 41559 40004 41604 40032
rect 36780 39992 36786 40004
rect 41598 39992 41604 40004
rect 41656 39992 41662 40044
rect 41782 40032 41788 40044
rect 41743 40004 41788 40032
rect 41782 39992 41788 40004
rect 41840 39992 41846 40044
rect 42797 40035 42855 40041
rect 42797 40001 42809 40035
rect 42843 40032 42855 40035
rect 43088 40032 43116 40072
rect 43162 40060 43168 40072
rect 43220 40060 43226 40112
rect 44082 40032 44088 40044
rect 42843 40004 43116 40032
rect 44043 40004 44088 40032
rect 42843 40001 42855 40004
rect 42797 39995 42855 40001
rect 44082 39992 44088 40004
rect 44140 39992 44146 40044
rect 45002 40041 45008 40044
rect 44996 39995 45008 40041
rect 45060 40032 45066 40044
rect 47762 40032 47768 40044
rect 45060 40004 45096 40032
rect 47723 40004 47768 40032
rect 45002 39992 45008 39995
rect 45060 39992 45066 40004
rect 47762 39992 47768 40004
rect 47820 39992 47826 40044
rect 35802 39964 35808 39976
rect 35268 39936 35480 39964
rect 35763 39936 35808 39964
rect 30745 39927 30803 39933
rect 35802 39924 35808 39936
rect 35860 39924 35866 39976
rect 38102 39924 38108 39976
rect 38160 39964 38166 39976
rect 38562 39964 38568 39976
rect 38160 39936 38568 39964
rect 38160 39924 38166 39936
rect 38562 39924 38568 39936
rect 38620 39964 38626 39976
rect 38657 39967 38715 39973
rect 38657 39964 38669 39967
rect 38620 39936 38669 39964
rect 38620 39924 38626 39936
rect 38657 39933 38669 39936
rect 38703 39933 38715 39967
rect 38657 39927 38715 39933
rect 41417 39967 41475 39973
rect 41417 39933 41429 39967
rect 41463 39964 41475 39967
rect 42613 39967 42671 39973
rect 42613 39964 42625 39967
rect 41463 39936 42625 39964
rect 41463 39933 41475 39936
rect 41417 39927 41475 39933
rect 42613 39933 42625 39936
rect 42659 39964 42671 39967
rect 43070 39964 43076 39976
rect 42659 39936 43076 39964
rect 42659 39933 42671 39936
rect 42613 39927 42671 39933
rect 43070 39924 43076 39936
rect 43128 39924 43134 39976
rect 43901 39967 43959 39973
rect 43901 39933 43913 39967
rect 43947 39964 43959 39967
rect 44174 39964 44180 39976
rect 43947 39936 44180 39964
rect 43947 39933 43959 39936
rect 43901 39927 43959 39933
rect 44174 39924 44180 39936
rect 44232 39924 44238 39976
rect 44726 39964 44732 39976
rect 44687 39936 44732 39964
rect 44726 39924 44732 39936
rect 44784 39924 44790 39976
rect 30374 39896 30380 39908
rect 29564 39868 30380 39896
rect 29564 39828 29592 39868
rect 30374 39856 30380 39868
rect 30432 39856 30438 39908
rect 35434 39856 35440 39908
rect 35492 39896 35498 39908
rect 36541 39899 36599 39905
rect 36541 39896 36553 39899
rect 35492 39868 36553 39896
rect 35492 39856 35498 39868
rect 36541 39865 36553 39868
rect 36587 39865 36599 39899
rect 36541 39859 36599 39865
rect 30466 39828 30472 39840
rect 27264 39800 29592 39828
rect 30427 39800 30472 39828
rect 30466 39788 30472 39800
rect 30524 39788 30530 39840
rect 35161 39831 35219 39837
rect 35161 39797 35173 39831
rect 35207 39828 35219 39831
rect 35710 39828 35716 39840
rect 35207 39800 35716 39828
rect 35207 39797 35219 39800
rect 35161 39791 35219 39797
rect 35710 39788 35716 39800
rect 35768 39788 35774 39840
rect 42794 39788 42800 39840
rect 42852 39828 42858 39840
rect 43165 39831 43223 39837
rect 43165 39828 43177 39831
rect 42852 39800 43177 39828
rect 42852 39788 42858 39800
rect 43165 39797 43177 39800
rect 43211 39797 43223 39831
rect 43165 39791 43223 39797
rect 44269 39831 44327 39837
rect 44269 39797 44281 39831
rect 44315 39828 44327 39831
rect 45370 39828 45376 39840
rect 44315 39800 45376 39828
rect 44315 39797 44327 39800
rect 44269 39791 44327 39797
rect 45370 39788 45376 39800
rect 45428 39788 45434 39840
rect 46474 39788 46480 39840
rect 46532 39828 46538 39840
rect 47213 39831 47271 39837
rect 47213 39828 47225 39831
rect 46532 39800 47225 39828
rect 46532 39788 46538 39800
rect 47213 39797 47225 39800
rect 47259 39797 47271 39831
rect 47854 39828 47860 39840
rect 47815 39800 47860 39828
rect 47213 39791 47271 39797
rect 47854 39788 47860 39800
rect 47912 39788 47918 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 23845 39627 23903 39633
rect 23845 39593 23857 39627
rect 23891 39624 23903 39627
rect 23934 39624 23940 39636
rect 23891 39596 23940 39624
rect 23891 39593 23903 39596
rect 23845 39587 23903 39593
rect 23934 39584 23940 39596
rect 23992 39584 23998 39636
rect 30006 39584 30012 39636
rect 30064 39624 30070 39636
rect 30101 39627 30159 39633
rect 30101 39624 30113 39627
rect 30064 39596 30113 39624
rect 30064 39584 30070 39596
rect 30101 39593 30113 39596
rect 30147 39593 30159 39627
rect 30101 39587 30159 39593
rect 32861 39627 32919 39633
rect 32861 39593 32873 39627
rect 32907 39624 32919 39627
rect 33226 39624 33232 39636
rect 32907 39596 33232 39624
rect 32907 39593 32919 39596
rect 32861 39587 32919 39593
rect 33226 39584 33232 39596
rect 33284 39584 33290 39636
rect 33962 39584 33968 39636
rect 34020 39624 34026 39636
rect 34241 39627 34299 39633
rect 34241 39624 34253 39627
rect 34020 39596 34253 39624
rect 34020 39584 34026 39596
rect 34241 39593 34253 39596
rect 34287 39593 34299 39627
rect 34241 39587 34299 39593
rect 35069 39627 35127 39633
rect 35069 39593 35081 39627
rect 35115 39593 35127 39627
rect 35434 39624 35440 39636
rect 35395 39596 35440 39624
rect 35069 39587 35127 39593
rect 24578 39516 24584 39568
rect 24636 39556 24642 39568
rect 35084 39556 35112 39587
rect 35434 39584 35440 39596
rect 35492 39584 35498 39636
rect 42337 39627 42395 39633
rect 42337 39593 42349 39627
rect 42383 39624 42395 39627
rect 42978 39624 42984 39636
rect 42383 39596 42984 39624
rect 42383 39593 42395 39596
rect 42337 39587 42395 39593
rect 42978 39584 42984 39596
rect 43036 39584 43042 39636
rect 45002 39584 45008 39636
rect 45060 39624 45066 39636
rect 45189 39627 45247 39633
rect 45189 39624 45201 39627
rect 45060 39596 45201 39624
rect 45060 39584 45066 39596
rect 45189 39593 45201 39596
rect 45235 39593 45247 39627
rect 45189 39587 45247 39593
rect 24636 39528 25544 39556
rect 24636 39516 24642 39528
rect 24949 39491 25007 39497
rect 24949 39488 24961 39491
rect 24044 39460 24961 39488
rect 24044 39429 24072 39460
rect 24949 39457 24961 39460
rect 24995 39457 25007 39491
rect 24949 39451 25007 39457
rect 24029 39423 24087 39429
rect 24029 39389 24041 39423
rect 24075 39389 24087 39423
rect 24029 39383 24087 39389
rect 24673 39423 24731 39429
rect 24673 39389 24685 39423
rect 24719 39389 24731 39423
rect 24673 39383 24731 39389
rect 24688 39284 24716 39383
rect 24762 39380 24768 39432
rect 24820 39420 24826 39432
rect 25516 39429 25544 39528
rect 33888 39528 35112 39556
rect 27433 39491 27491 39497
rect 27433 39457 27445 39491
rect 27479 39488 27491 39491
rect 28258 39488 28264 39500
rect 27479 39460 28264 39488
rect 27479 39457 27491 39460
rect 27433 39451 27491 39457
rect 28258 39448 28264 39460
rect 28316 39448 28322 39500
rect 30098 39488 30104 39500
rect 28460 39460 30104 39488
rect 25501 39423 25559 39429
rect 24820 39392 24865 39420
rect 24820 39380 24826 39392
rect 25501 39389 25513 39423
rect 25547 39389 25559 39423
rect 25501 39383 25559 39389
rect 27617 39423 27675 39429
rect 27617 39389 27629 39423
rect 27663 39420 27675 39423
rect 28166 39420 28172 39432
rect 27663 39392 28172 39420
rect 27663 39389 27675 39392
rect 27617 39383 27675 39389
rect 28166 39380 28172 39392
rect 28224 39380 28230 39432
rect 28460 39429 28488 39460
rect 30098 39448 30104 39460
rect 30156 39448 30162 39500
rect 28445 39423 28503 39429
rect 28445 39389 28457 39423
rect 28491 39389 28503 39423
rect 28626 39420 28632 39432
rect 28587 39392 28632 39420
rect 28445 39383 28503 39389
rect 28626 39380 28632 39392
rect 28684 39380 28690 39432
rect 28902 39420 28908 39432
rect 28863 39392 28908 39420
rect 28902 39380 28908 39392
rect 28960 39380 28966 39432
rect 29730 39420 29736 39432
rect 29691 39392 29736 39420
rect 29730 39380 29736 39392
rect 29788 39380 29794 39432
rect 29917 39423 29975 39429
rect 29917 39389 29929 39423
rect 29963 39420 29975 39423
rect 30374 39420 30380 39432
rect 29963 39392 30380 39420
rect 29963 39389 29975 39392
rect 29917 39383 29975 39389
rect 30374 39380 30380 39392
rect 30432 39420 30438 39432
rect 31294 39420 31300 39432
rect 30432 39392 31300 39420
rect 30432 39380 30438 39392
rect 31294 39380 31300 39392
rect 31352 39380 31358 39432
rect 31478 39380 31484 39432
rect 31536 39420 31542 39432
rect 31941 39423 31999 39429
rect 31941 39420 31953 39423
rect 31536 39392 31953 39420
rect 31536 39380 31542 39392
rect 31941 39389 31953 39392
rect 31987 39389 31999 39423
rect 31941 39383 31999 39389
rect 25768 39355 25826 39361
rect 25768 39321 25780 39355
rect 25814 39352 25826 39355
rect 26418 39352 26424 39364
rect 25814 39324 26424 39352
rect 25814 39321 25826 39324
rect 25768 39315 25826 39321
rect 26418 39312 26424 39324
rect 26476 39312 26482 39364
rect 28534 39352 28540 39364
rect 28495 39324 28540 39352
rect 28534 39312 28540 39324
rect 28592 39312 28598 39364
rect 28767 39355 28825 39361
rect 28767 39321 28779 39355
rect 28813 39352 28825 39355
rect 30466 39352 30472 39364
rect 28813 39324 30472 39352
rect 28813 39321 28825 39324
rect 28767 39315 28825 39321
rect 30466 39312 30472 39324
rect 30524 39312 30530 39364
rect 31956 39352 31984 39383
rect 32030 39380 32036 39432
rect 32088 39420 32094 39432
rect 32125 39423 32183 39429
rect 32125 39420 32137 39423
rect 32088 39392 32137 39420
rect 32088 39380 32094 39392
rect 32125 39389 32137 39392
rect 32171 39389 32183 39423
rect 32125 39383 32183 39389
rect 32309 39423 32367 39429
rect 32309 39389 32321 39423
rect 32355 39420 32367 39423
rect 33045 39423 33103 39429
rect 33045 39420 33057 39423
rect 32355 39392 33057 39420
rect 32355 39389 32367 39392
rect 32309 39383 32367 39389
rect 33045 39389 33057 39392
rect 33091 39389 33103 39423
rect 33045 39383 33103 39389
rect 33888 39352 33916 39528
rect 35526 39488 35532 39500
rect 35084 39460 35532 39488
rect 33965 39423 34023 39429
rect 33965 39389 33977 39423
rect 34011 39389 34023 39423
rect 33965 39383 34023 39389
rect 31956 39324 33916 39352
rect 33980 39352 34008 39383
rect 34054 39380 34060 39432
rect 34112 39420 34118 39432
rect 35084 39429 35112 39460
rect 35526 39448 35532 39460
rect 35584 39448 35590 39500
rect 46474 39488 46480 39500
rect 46435 39460 46480 39488
rect 46474 39448 46480 39460
rect 46532 39448 46538 39500
rect 46661 39491 46719 39497
rect 46661 39457 46673 39491
rect 46707 39488 46719 39491
rect 47854 39488 47860 39500
rect 46707 39460 47860 39488
rect 46707 39457 46719 39460
rect 46661 39451 46719 39457
rect 47854 39448 47860 39460
rect 47912 39448 47918 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 35069 39423 35127 39429
rect 34112 39392 34157 39420
rect 34112 39380 34118 39392
rect 35069 39389 35081 39423
rect 35115 39389 35127 39423
rect 35069 39383 35127 39389
rect 35161 39423 35219 39429
rect 35161 39389 35173 39423
rect 35207 39389 35219 39423
rect 38102 39420 38108 39432
rect 38063 39392 38108 39420
rect 35161 39383 35219 39389
rect 34514 39352 34520 39364
rect 33980 39324 34520 39352
rect 34514 39312 34520 39324
rect 34572 39352 34578 39364
rect 35176 39352 35204 39383
rect 38102 39380 38108 39392
rect 38160 39380 38166 39432
rect 38372 39423 38430 39429
rect 38372 39389 38384 39423
rect 38418 39420 38430 39423
rect 39666 39420 39672 39432
rect 38418 39392 39672 39420
rect 38418 39389 38430 39392
rect 38372 39383 38430 39389
rect 39666 39380 39672 39392
rect 39724 39380 39730 39432
rect 42518 39420 42524 39432
rect 42479 39392 42524 39420
rect 42518 39380 42524 39392
rect 42576 39380 42582 39432
rect 45370 39420 45376 39432
rect 45331 39392 45376 39420
rect 45370 39380 45376 39392
rect 45428 39380 45434 39432
rect 34572 39324 35204 39352
rect 36725 39355 36783 39361
rect 34572 39312 34578 39324
rect 36725 39321 36737 39355
rect 36771 39352 36783 39355
rect 37550 39352 37556 39364
rect 36771 39324 37556 39352
rect 36771 39321 36783 39324
rect 36725 39315 36783 39321
rect 37550 39312 37556 39324
rect 37608 39312 37614 39364
rect 25590 39284 25596 39296
rect 24688 39256 25596 39284
rect 25590 39244 25596 39256
rect 25648 39244 25654 39296
rect 25682 39244 25688 39296
rect 25740 39284 25746 39296
rect 26881 39287 26939 39293
rect 26881 39284 26893 39287
rect 25740 39256 26893 39284
rect 25740 39244 25746 39256
rect 26881 39253 26893 39256
rect 26927 39253 26939 39287
rect 27798 39284 27804 39296
rect 27759 39256 27804 39284
rect 26881 39247 26939 39253
rect 27798 39244 27804 39256
rect 27856 39244 27862 39296
rect 28261 39287 28319 39293
rect 28261 39253 28273 39287
rect 28307 39284 28319 39287
rect 28350 39284 28356 39296
rect 28307 39256 28356 39284
rect 28307 39253 28319 39256
rect 28261 39247 28319 39253
rect 28350 39244 28356 39256
rect 28408 39244 28414 39296
rect 34054 39244 34060 39296
rect 34112 39284 34118 39296
rect 36817 39287 36875 39293
rect 36817 39284 36829 39287
rect 34112 39256 36829 39284
rect 34112 39244 34118 39256
rect 36817 39253 36829 39256
rect 36863 39253 36875 39287
rect 36817 39247 36875 39253
rect 38654 39244 38660 39296
rect 38712 39284 38718 39296
rect 39485 39287 39543 39293
rect 39485 39284 39497 39287
rect 38712 39256 39497 39284
rect 38712 39244 38718 39256
rect 39485 39253 39497 39256
rect 39531 39253 39543 39287
rect 39485 39247 39543 39253
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 25682 39080 25688 39092
rect 25643 39052 25688 39080
rect 25682 39040 25688 39052
rect 25740 39040 25746 39092
rect 25774 39040 25780 39092
rect 25832 39080 25838 39092
rect 26418 39080 26424 39092
rect 25832 39052 25877 39080
rect 26379 39052 26424 39080
rect 25832 39040 25838 39052
rect 26418 39040 26424 39052
rect 26476 39040 26482 39092
rect 29457 39083 29515 39089
rect 29457 39049 29469 39083
rect 29503 39080 29515 39083
rect 29730 39080 29736 39092
rect 29503 39052 29736 39080
rect 29503 39049 29515 39052
rect 29457 39043 29515 39049
rect 29730 39040 29736 39052
rect 29788 39040 29794 39092
rect 32493 39083 32551 39089
rect 32493 39049 32505 39083
rect 32539 39080 32551 39083
rect 32539 39052 33180 39080
rect 32539 39049 32551 39052
rect 32493 39043 32551 39049
rect 25038 38972 25044 39024
rect 25096 39012 25102 39024
rect 25409 39015 25467 39021
rect 25409 39012 25421 39015
rect 25096 38984 25421 39012
rect 25096 38972 25102 38984
rect 25409 38981 25421 38984
rect 25455 38981 25467 39015
rect 25590 39012 25596 39024
rect 25551 38984 25596 39012
rect 25409 38975 25467 38981
rect 25590 38972 25596 38984
rect 25648 38972 25654 39024
rect 28344 39015 28402 39021
rect 28344 38981 28356 39015
rect 28390 39012 28402 39015
rect 28534 39012 28540 39024
rect 28390 38984 28540 39012
rect 28390 38981 28402 38984
rect 28344 38975 28402 38981
rect 28534 38972 28540 38984
rect 28592 38972 28598 39024
rect 28902 38972 28908 39024
rect 28960 39012 28966 39024
rect 28960 38984 32444 39012
rect 28960 38972 28966 38984
rect 26602 38944 26608 38956
rect 26563 38916 26608 38944
rect 26602 38904 26608 38916
rect 26660 38904 26666 38956
rect 28074 38944 28080 38956
rect 28035 38916 28080 38944
rect 28074 38904 28080 38916
rect 28132 38904 28138 38956
rect 31202 38944 31208 38956
rect 31163 38916 31208 38944
rect 31202 38904 31208 38916
rect 31260 38904 31266 38956
rect 32030 38904 32036 38956
rect 32088 38944 32094 38956
rect 32309 38947 32367 38953
rect 32309 38944 32321 38947
rect 32088 38916 32321 38944
rect 32088 38904 32094 38916
rect 32309 38913 32321 38916
rect 32355 38913 32367 38947
rect 32416 38944 32444 38984
rect 33152 38953 33180 39052
rect 36722 39040 36728 39092
rect 36780 39080 36786 39092
rect 36817 39083 36875 39089
rect 36817 39080 36829 39083
rect 36780 39052 36829 39080
rect 36780 39040 36786 39052
rect 36817 39049 36829 39052
rect 36863 39049 36875 39083
rect 36817 39043 36875 39049
rect 39301 39083 39359 39089
rect 39301 39049 39313 39083
rect 39347 39080 39359 39083
rect 40218 39080 40224 39092
rect 39347 39052 40224 39080
rect 39347 39049 39359 39052
rect 39301 39043 39359 39049
rect 40218 39040 40224 39052
rect 40276 39040 40282 39092
rect 44637 39083 44695 39089
rect 44637 39080 44649 39083
rect 43548 39052 44649 39080
rect 35710 39021 35716 39024
rect 35704 39012 35716 39021
rect 35671 38984 35716 39012
rect 35704 38975 35716 38984
rect 35710 38972 35716 38975
rect 35768 38972 35774 39024
rect 43254 38972 43260 39024
rect 43312 39012 43318 39024
rect 43548 39021 43576 39052
rect 44637 39049 44649 39052
rect 44683 39049 44695 39083
rect 44637 39043 44695 39049
rect 45189 39083 45247 39089
rect 45189 39049 45201 39083
rect 45235 39049 45247 39083
rect 45189 39043 45247 39049
rect 43349 39015 43407 39021
rect 43349 39012 43361 39015
rect 43312 38984 43361 39012
rect 43312 38972 43318 38984
rect 43349 38981 43361 38984
rect 43395 38981 43407 39015
rect 43349 38975 43407 38981
rect 43533 39015 43591 39021
rect 43533 38981 43545 39015
rect 43579 38981 43591 39015
rect 45204 39012 45232 39043
rect 46078 39015 46136 39021
rect 46078 39012 46090 39015
rect 45204 38984 46090 39012
rect 43533 38975 43591 38981
rect 46078 38981 46090 38984
rect 46124 38981 46136 39015
rect 46078 38975 46136 38981
rect 33137 38947 33195 38953
rect 32416 38916 32996 38944
rect 32309 38907 32367 38913
rect 32968 38808 32996 38916
rect 33137 38913 33149 38947
rect 33183 38944 33195 38947
rect 37550 38944 37556 38956
rect 33183 38916 37556 38944
rect 33183 38913 33195 38916
rect 33137 38907 33195 38913
rect 37550 38904 37556 38916
rect 37608 38944 37614 38956
rect 37737 38947 37795 38953
rect 37737 38944 37749 38947
rect 37608 38916 37749 38944
rect 37608 38904 37614 38916
rect 37737 38913 37749 38916
rect 37783 38944 37795 38947
rect 39022 38944 39028 38956
rect 37783 38916 39028 38944
rect 37783 38913 37795 38916
rect 37737 38907 37795 38913
rect 39022 38904 39028 38916
rect 39080 38944 39086 38956
rect 39209 38947 39267 38953
rect 39209 38944 39221 38947
rect 39080 38916 39221 38944
rect 39080 38904 39086 38916
rect 39209 38913 39221 38916
rect 39255 38913 39267 38947
rect 44174 38944 44180 38956
rect 44087 38916 44180 38944
rect 39209 38907 39267 38913
rect 44174 38904 44180 38916
rect 44232 38904 44238 38956
rect 44450 38944 44456 38956
rect 44411 38916 44456 38944
rect 44450 38904 44456 38916
rect 44508 38904 44514 38956
rect 45373 38947 45431 38953
rect 45373 38913 45385 38947
rect 45419 38944 45431 38947
rect 45554 38944 45560 38956
rect 45419 38916 45560 38944
rect 45419 38913 45431 38916
rect 45373 38907 45431 38913
rect 45554 38904 45560 38916
rect 45612 38904 45618 38956
rect 33042 38836 33048 38888
rect 33100 38876 33106 38888
rect 35437 38879 35495 38885
rect 35437 38876 35449 38879
rect 33100 38848 35449 38876
rect 33100 38836 33106 38848
rect 35437 38845 35449 38848
rect 35483 38845 35495 38879
rect 35437 38839 35495 38845
rect 37921 38879 37979 38885
rect 37921 38845 37933 38879
rect 37967 38876 37979 38879
rect 43530 38876 43536 38888
rect 37967 38848 43536 38876
rect 37967 38845 37979 38848
rect 37921 38839 37979 38845
rect 34606 38808 34612 38820
rect 32416 38780 32904 38808
rect 32968 38780 34612 38808
rect 25958 38740 25964 38752
rect 25919 38712 25964 38740
rect 25958 38700 25964 38712
rect 26016 38700 26022 38752
rect 31021 38743 31079 38749
rect 31021 38709 31033 38743
rect 31067 38740 31079 38743
rect 31110 38740 31116 38752
rect 31067 38712 31116 38740
rect 31067 38709 31079 38712
rect 31021 38703 31079 38709
rect 31110 38700 31116 38712
rect 31168 38700 31174 38752
rect 31294 38700 31300 38752
rect 31352 38740 31358 38752
rect 32416 38740 32444 38780
rect 32876 38752 32904 38780
rect 34606 38768 34612 38780
rect 34664 38768 34670 38820
rect 31352 38712 32444 38740
rect 31352 38700 31358 38712
rect 32858 38700 32864 38752
rect 32916 38740 32922 38752
rect 33229 38743 33287 38749
rect 33229 38740 33241 38743
rect 32916 38712 33241 38740
rect 32916 38700 32922 38712
rect 33229 38709 33241 38712
rect 33275 38709 33287 38743
rect 34624 38740 34652 38768
rect 35802 38740 35808 38752
rect 34624 38712 35808 38740
rect 33229 38703 33287 38709
rect 35802 38700 35808 38712
rect 35860 38740 35866 38752
rect 37936 38740 37964 38839
rect 43530 38836 43536 38848
rect 43588 38836 43594 38888
rect 44192 38808 44220 38904
rect 44358 38876 44364 38888
rect 44271 38848 44364 38876
rect 44358 38836 44364 38848
rect 44416 38876 44422 38888
rect 45278 38876 45284 38888
rect 44416 38848 45284 38876
rect 44416 38836 44422 38848
rect 45278 38836 45284 38848
rect 45336 38836 45342 38888
rect 45462 38836 45468 38888
rect 45520 38876 45526 38888
rect 45833 38879 45891 38885
rect 45833 38876 45845 38879
rect 45520 38848 45845 38876
rect 45520 38836 45526 38848
rect 45833 38845 45845 38848
rect 45879 38845 45891 38879
rect 45833 38839 45891 38845
rect 44192 38780 44404 38808
rect 43714 38740 43720 38752
rect 35860 38712 37964 38740
rect 43675 38712 43720 38740
rect 35860 38700 35866 38712
rect 43714 38700 43720 38712
rect 43772 38700 43778 38752
rect 44266 38740 44272 38752
rect 44227 38712 44272 38740
rect 44266 38700 44272 38712
rect 44324 38700 44330 38752
rect 44376 38740 44404 38780
rect 44542 38740 44548 38752
rect 44376 38712 44548 38740
rect 44542 38700 44548 38712
rect 44600 38740 44606 38752
rect 47213 38743 47271 38749
rect 47213 38740 47225 38743
rect 44600 38712 47225 38740
rect 44600 38700 44606 38712
rect 47213 38709 47225 38712
rect 47259 38709 47271 38743
rect 47946 38740 47952 38752
rect 47907 38712 47952 38740
rect 47213 38703 47271 38709
rect 47946 38700 47952 38712
rect 48004 38700 48010 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 25590 38536 25596 38548
rect 25551 38508 25596 38536
rect 25590 38496 25596 38508
rect 25648 38496 25654 38548
rect 28534 38536 28540 38548
rect 28495 38508 28540 38536
rect 28534 38496 28540 38508
rect 28592 38496 28598 38548
rect 32122 38536 32128 38548
rect 30852 38508 32128 38536
rect 25682 38400 25688 38412
rect 25643 38372 25688 38400
rect 25682 38360 25688 38372
rect 25740 38360 25746 38412
rect 30852 38409 30880 38508
rect 32122 38496 32128 38508
rect 32180 38496 32186 38548
rect 40034 38536 40040 38548
rect 39947 38508 40040 38536
rect 40034 38496 40040 38508
rect 40092 38536 40098 38548
rect 45554 38536 45560 38548
rect 40092 38508 43208 38536
rect 45515 38508 45560 38536
rect 40092 38496 40098 38508
rect 32217 38471 32275 38477
rect 32217 38437 32229 38471
rect 32263 38468 32275 38471
rect 32263 38440 32720 38468
rect 32263 38437 32275 38440
rect 32217 38431 32275 38437
rect 32692 38409 32720 38440
rect 30837 38403 30895 38409
rect 30837 38369 30849 38403
rect 30883 38369 30895 38403
rect 30837 38363 30895 38369
rect 32677 38403 32735 38409
rect 32677 38369 32689 38403
rect 32723 38400 32735 38403
rect 33410 38400 33416 38412
rect 32723 38372 33416 38400
rect 32723 38369 32735 38372
rect 32677 38363 32735 38369
rect 33410 38360 33416 38372
rect 33468 38360 33474 38412
rect 36722 38360 36728 38412
rect 36780 38400 36786 38412
rect 36909 38403 36967 38409
rect 36909 38400 36921 38403
rect 36780 38372 36921 38400
rect 36780 38360 36786 38372
rect 36909 38369 36921 38372
rect 36955 38400 36967 38403
rect 37182 38400 37188 38412
rect 36955 38372 37188 38400
rect 36955 38369 36967 38372
rect 36909 38363 36967 38369
rect 37182 38360 37188 38372
rect 37240 38360 37246 38412
rect 43070 38400 43076 38412
rect 42628 38372 43076 38400
rect 24762 38332 24768 38344
rect 24723 38304 24768 38332
rect 24762 38292 24768 38304
rect 24820 38292 24826 38344
rect 25038 38292 25044 38344
rect 25096 38332 25102 38344
rect 25777 38335 25835 38341
rect 25777 38332 25789 38335
rect 25096 38304 25789 38332
rect 25096 38292 25102 38304
rect 25777 38301 25789 38304
rect 25823 38301 25835 38335
rect 25777 38295 25835 38301
rect 27798 38292 27804 38344
rect 27856 38332 27862 38344
rect 31110 38341 31116 38344
rect 28721 38335 28779 38341
rect 28721 38332 28733 38335
rect 27856 38304 28733 38332
rect 27856 38292 27862 38304
rect 28721 38301 28733 38304
rect 28767 38301 28779 38335
rect 31104 38332 31116 38341
rect 31071 38304 31116 38332
rect 28721 38295 28779 38301
rect 31104 38295 31116 38304
rect 31110 38292 31116 38295
rect 31168 38292 31174 38344
rect 32858 38332 32864 38344
rect 32819 38304 32864 38332
rect 32858 38292 32864 38304
rect 32916 38292 32922 38344
rect 33045 38335 33103 38341
rect 33045 38301 33057 38335
rect 33091 38332 33103 38335
rect 33689 38335 33747 38341
rect 33689 38332 33701 38335
rect 33091 38304 33701 38332
rect 33091 38301 33103 38304
rect 33045 38295 33103 38301
rect 33689 38301 33701 38304
rect 33735 38301 33747 38335
rect 37090 38332 37096 38344
rect 37003 38304 37096 38332
rect 33689 38295 33747 38301
rect 37090 38292 37096 38304
rect 37148 38332 37154 38344
rect 38746 38332 38752 38344
rect 37148 38304 38752 38332
rect 37148 38292 37154 38304
rect 38746 38292 38752 38304
rect 38804 38292 38810 38344
rect 38933 38335 38991 38341
rect 38933 38301 38945 38335
rect 38979 38301 38991 38335
rect 38933 38295 38991 38301
rect 25501 38267 25559 38273
rect 25501 38233 25513 38267
rect 25547 38264 25559 38267
rect 25682 38264 25688 38276
rect 25547 38236 25688 38264
rect 25547 38233 25559 38236
rect 25501 38227 25559 38233
rect 25682 38224 25688 38236
rect 25740 38224 25746 38276
rect 38948 38264 38976 38295
rect 39022 38292 39028 38344
rect 39080 38332 39086 38344
rect 39209 38335 39267 38341
rect 39080 38304 39125 38332
rect 39080 38292 39086 38304
rect 39209 38301 39221 38335
rect 39255 38332 39267 38335
rect 40221 38335 40279 38341
rect 40221 38332 40233 38335
rect 39255 38304 40233 38332
rect 39255 38301 39267 38304
rect 39209 38295 39267 38301
rect 40221 38301 40233 38304
rect 40267 38301 40279 38335
rect 40221 38295 40279 38301
rect 40681 38335 40739 38341
rect 40681 38301 40693 38335
rect 40727 38332 40739 38335
rect 42628 38332 42656 38372
rect 43070 38360 43076 38372
rect 43128 38360 43134 38412
rect 40727 38304 42656 38332
rect 42705 38335 42763 38341
rect 40727 38301 40739 38304
rect 40681 38295 40739 38301
rect 42705 38301 42717 38335
rect 42751 38301 42763 38335
rect 42705 38295 42763 38301
rect 40948 38267 41006 38273
rect 38948 38236 39988 38264
rect 39960 38208 39988 38236
rect 40948 38233 40960 38267
rect 40994 38264 41006 38267
rect 42521 38267 42579 38273
rect 42521 38264 42533 38267
rect 40994 38236 42533 38264
rect 40994 38233 41006 38236
rect 40948 38227 41006 38233
rect 42521 38233 42533 38236
rect 42567 38233 42579 38267
rect 42521 38227 42579 38233
rect 23842 38156 23848 38208
rect 23900 38196 23906 38208
rect 24581 38199 24639 38205
rect 24581 38196 24593 38199
rect 23900 38168 24593 38196
rect 23900 38156 23906 38168
rect 24581 38165 24593 38168
rect 24627 38165 24639 38199
rect 24581 38159 24639 38165
rect 25961 38199 26019 38205
rect 25961 38165 25973 38199
rect 26007 38196 26019 38199
rect 26234 38196 26240 38208
rect 26007 38168 26240 38196
rect 26007 38165 26019 38168
rect 25961 38159 26019 38165
rect 26234 38156 26240 38168
rect 26292 38156 26298 38208
rect 33502 38196 33508 38208
rect 33463 38168 33508 38196
rect 33502 38156 33508 38168
rect 33560 38156 33566 38208
rect 36906 38156 36912 38208
rect 36964 38196 36970 38208
rect 37277 38199 37335 38205
rect 37277 38196 37289 38199
rect 36964 38168 37289 38196
rect 36964 38156 36970 38168
rect 37277 38165 37289 38168
rect 37323 38165 37335 38199
rect 37277 38159 37335 38165
rect 39942 38156 39948 38208
rect 40000 38196 40006 38208
rect 42061 38199 42119 38205
rect 42061 38196 42073 38199
rect 40000 38168 42073 38196
rect 40000 38156 40006 38168
rect 42061 38165 42073 38168
rect 42107 38165 42119 38199
rect 42720 38196 42748 38295
rect 42794 38292 42800 38344
rect 42852 38332 42858 38344
rect 43180 38341 43208 38508
rect 45554 38496 45560 38508
rect 45612 38496 45618 38548
rect 44085 38471 44143 38477
rect 44085 38437 44097 38471
rect 44131 38468 44143 38471
rect 44450 38468 44456 38480
rect 44131 38440 44456 38468
rect 44131 38437 44143 38440
rect 44085 38431 44143 38437
rect 44450 38428 44456 38440
rect 44508 38468 44514 38480
rect 45094 38468 45100 38480
rect 44508 38440 45100 38468
rect 44508 38428 44514 38440
rect 45094 38428 45100 38440
rect 45152 38428 45158 38480
rect 43346 38360 43352 38412
rect 43404 38400 43410 38412
rect 44726 38400 44732 38412
rect 43404 38372 44732 38400
rect 43404 38360 43410 38372
rect 44726 38360 44732 38372
rect 44784 38400 44790 38412
rect 45462 38400 45468 38412
rect 44784 38372 45468 38400
rect 44784 38360 44790 38372
rect 45462 38360 45468 38372
rect 45520 38360 45526 38412
rect 48038 38400 48044 38412
rect 47999 38372 48044 38400
rect 48038 38360 48044 38372
rect 48096 38360 48102 38412
rect 43165 38335 43223 38341
rect 42852 38304 42897 38332
rect 42852 38292 42858 38304
rect 43165 38301 43177 38335
rect 43211 38301 43223 38335
rect 44266 38332 44272 38344
rect 44227 38304 44272 38332
rect 43165 38295 43223 38301
rect 44266 38292 44272 38304
rect 44324 38292 44330 38344
rect 44358 38292 44364 38344
rect 44416 38332 44422 38344
rect 44416 38304 44461 38332
rect 44416 38292 44422 38304
rect 45094 38292 45100 38344
rect 45152 38332 45158 38344
rect 45189 38335 45247 38341
rect 45189 38332 45201 38335
rect 45152 38304 45201 38332
rect 45152 38292 45158 38304
rect 45189 38301 45201 38304
rect 45235 38301 45247 38335
rect 45370 38332 45376 38344
rect 45331 38304 45376 38332
rect 45189 38295 45247 38301
rect 45370 38292 45376 38304
rect 45428 38292 45434 38344
rect 46106 38292 46112 38344
rect 46164 38332 46170 38344
rect 46477 38335 46535 38341
rect 46477 38332 46489 38335
rect 46164 38304 46489 38332
rect 46164 38292 46170 38304
rect 46477 38301 46489 38304
rect 46523 38301 46535 38335
rect 46477 38295 46535 38301
rect 42886 38264 42892 38276
rect 42847 38236 42892 38264
rect 42886 38224 42892 38236
rect 42944 38224 42950 38276
rect 43027 38267 43085 38273
rect 43027 38233 43039 38267
rect 43073 38264 43085 38267
rect 43714 38264 43720 38276
rect 43073 38236 43720 38264
rect 43073 38233 43085 38236
rect 43027 38227 43085 38233
rect 43714 38224 43720 38236
rect 43772 38224 43778 38276
rect 44637 38267 44695 38273
rect 44637 38264 44649 38267
rect 44192 38236 44649 38264
rect 44192 38196 44220 38236
rect 44637 38233 44649 38236
rect 44683 38233 44695 38267
rect 44637 38227 44695 38233
rect 46661 38267 46719 38273
rect 46661 38233 46673 38267
rect 46707 38264 46719 38267
rect 46842 38264 46848 38276
rect 46707 38236 46848 38264
rect 46707 38233 46719 38236
rect 46661 38227 46719 38233
rect 46842 38224 46848 38236
rect 46900 38224 46906 38276
rect 42720 38168 44220 38196
rect 44453 38199 44511 38205
rect 42061 38159 42119 38165
rect 44453 38165 44465 38199
rect 44499 38196 44511 38199
rect 44542 38196 44548 38208
rect 44499 38168 44548 38196
rect 44499 38165 44511 38168
rect 44453 38159 44511 38165
rect 44542 38156 44548 38168
rect 44600 38156 44606 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 24949 37995 25007 38001
rect 24949 37961 24961 37995
rect 24995 37992 25007 37995
rect 25590 37992 25596 38004
rect 24995 37964 25596 37992
rect 24995 37961 25007 37964
rect 24949 37955 25007 37961
rect 25590 37952 25596 37964
rect 25648 37952 25654 38004
rect 29454 37992 29460 38004
rect 29367 37964 29460 37992
rect 29454 37952 29460 37964
rect 29512 37992 29518 38004
rect 30926 37992 30932 38004
rect 29512 37964 30932 37992
rect 29512 37952 29518 37964
rect 30926 37952 30932 37964
rect 30984 37952 30990 38004
rect 31202 37952 31208 38004
rect 31260 37992 31266 38004
rect 31389 37995 31447 38001
rect 31389 37992 31401 37995
rect 31260 37964 31401 37992
rect 31260 37952 31266 37964
rect 31389 37961 31401 37964
rect 31435 37961 31447 37995
rect 31389 37955 31447 37961
rect 36725 37995 36783 38001
rect 36725 37961 36737 37995
rect 36771 37992 36783 37995
rect 43073 37995 43131 38001
rect 36771 37964 37596 37992
rect 36771 37961 36783 37964
rect 36725 37955 36783 37961
rect 23842 37933 23848 37936
rect 23836 37924 23848 37933
rect 23803 37896 23848 37924
rect 23836 37887 23848 37896
rect 23842 37884 23848 37887
rect 23900 37884 23906 37936
rect 32852 37927 32910 37933
rect 32852 37893 32864 37927
rect 32898 37924 32910 37927
rect 33502 37924 33508 37936
rect 32898 37896 33508 37924
rect 32898 37893 32910 37896
rect 32852 37887 32910 37893
rect 33502 37884 33508 37896
rect 33560 37884 33566 37936
rect 24578 37856 24584 37868
rect 23584 37828 24584 37856
rect 23584 37797 23612 37828
rect 24578 37816 24584 37828
rect 24636 37816 24642 37868
rect 28074 37856 28080 37868
rect 28035 37828 28080 37856
rect 28074 37816 28080 37828
rect 28132 37816 28138 37868
rect 28350 37865 28356 37868
rect 28344 37856 28356 37865
rect 28311 37828 28356 37856
rect 28344 37819 28356 37828
rect 28350 37816 28356 37819
rect 28408 37816 28414 37868
rect 31202 37856 31208 37868
rect 31163 37828 31208 37856
rect 31202 37816 31208 37828
rect 31260 37816 31266 37868
rect 32122 37816 32128 37868
rect 32180 37856 32186 37868
rect 32585 37859 32643 37865
rect 32585 37856 32597 37859
rect 32180 37828 32597 37856
rect 32180 37816 32186 37828
rect 32585 37825 32597 37828
rect 32631 37825 32643 37859
rect 36906 37856 36912 37868
rect 36867 37828 36912 37856
rect 32585 37819 32643 37825
rect 36906 37816 36912 37828
rect 36964 37816 36970 37868
rect 37568 37856 37596 37964
rect 43073 37961 43085 37995
rect 43119 37961 43131 37995
rect 45094 37992 45100 38004
rect 45055 37964 45100 37992
rect 43073 37955 43131 37961
rect 39936 37927 39994 37933
rect 39936 37893 39948 37927
rect 39982 37924 39994 37927
rect 40034 37924 40040 37936
rect 39982 37896 40040 37924
rect 39982 37893 39994 37896
rect 39936 37887 39994 37893
rect 40034 37884 40040 37896
rect 40092 37884 40098 37936
rect 43088 37924 43116 37955
rect 45094 37952 45100 37964
rect 45152 37952 45158 38004
rect 46106 37992 46112 38004
rect 46067 37964 46112 37992
rect 46106 37952 46112 37964
rect 46164 37952 46170 38004
rect 46842 37992 46848 38004
rect 46803 37964 46848 37992
rect 46842 37952 46848 37964
rect 46900 37952 46906 38004
rect 43962 37927 44020 37933
rect 43962 37924 43974 37927
rect 43088 37896 43974 37924
rect 43962 37893 43974 37896
rect 44008 37893 44020 37927
rect 43962 37887 44020 37893
rect 37717 37859 37775 37865
rect 37717 37856 37729 37859
rect 37568 37828 37729 37856
rect 37717 37825 37729 37828
rect 37763 37825 37775 37859
rect 39669 37859 39727 37865
rect 39669 37856 39681 37859
rect 37717 37819 37775 37825
rect 38488 37828 39681 37856
rect 23569 37791 23627 37797
rect 23569 37757 23581 37791
rect 23615 37757 23627 37791
rect 31018 37788 31024 37800
rect 30979 37760 31024 37788
rect 23569 37751 23627 37757
rect 31018 37748 31024 37760
rect 31076 37748 31082 37800
rect 37458 37788 37464 37800
rect 37419 37760 37464 37788
rect 37458 37748 37464 37760
rect 37516 37748 37522 37800
rect 33962 37652 33968 37664
rect 33923 37624 33968 37652
rect 33962 37612 33968 37624
rect 34020 37612 34026 37664
rect 37458 37612 37464 37664
rect 37516 37652 37522 37664
rect 38102 37652 38108 37664
rect 37516 37624 38108 37652
rect 37516 37612 37522 37624
rect 38102 37612 38108 37624
rect 38160 37652 38166 37664
rect 38488 37652 38516 37828
rect 39669 37825 39681 37828
rect 39715 37825 39727 37859
rect 39669 37819 39727 37825
rect 43257 37859 43315 37865
rect 43257 37825 43269 37859
rect 43303 37856 43315 37859
rect 44266 37856 44272 37868
rect 43303 37828 44272 37856
rect 43303 37825 43315 37828
rect 43257 37819 43315 37825
rect 44266 37816 44272 37828
rect 44324 37816 44330 37868
rect 46290 37856 46296 37868
rect 46251 37828 46296 37856
rect 46290 37816 46296 37828
rect 46348 37816 46354 37868
rect 46750 37856 46756 37868
rect 46711 37828 46756 37856
rect 46750 37816 46756 37828
rect 46808 37816 46814 37868
rect 47302 37816 47308 37868
rect 47360 37856 47366 37868
rect 47670 37856 47676 37868
rect 47360 37828 47676 37856
rect 47360 37816 47366 37828
rect 47670 37816 47676 37828
rect 47728 37856 47734 37868
rect 47765 37859 47823 37865
rect 47765 37856 47777 37859
rect 47728 37828 47777 37856
rect 47728 37816 47734 37828
rect 47765 37825 47777 37828
rect 47811 37825 47823 37859
rect 47765 37819 47823 37825
rect 43070 37748 43076 37800
rect 43128 37788 43134 37800
rect 43346 37788 43352 37800
rect 43128 37760 43352 37788
rect 43128 37748 43134 37760
rect 43346 37748 43352 37760
rect 43404 37788 43410 37800
rect 43717 37791 43775 37797
rect 43717 37788 43729 37791
rect 43404 37760 43729 37788
rect 43404 37748 43410 37760
rect 43717 37757 43729 37760
rect 43763 37757 43775 37791
rect 43717 37751 43775 37757
rect 38160 37624 38516 37652
rect 38841 37655 38899 37661
rect 38160 37612 38166 37624
rect 38841 37621 38853 37655
rect 38887 37652 38899 37655
rect 40310 37652 40316 37664
rect 38887 37624 40316 37652
rect 38887 37621 38899 37624
rect 38841 37615 38899 37621
rect 40310 37612 40316 37624
rect 40368 37612 40374 37664
rect 41046 37652 41052 37664
rect 41007 37624 41052 37652
rect 41046 37612 41052 37624
rect 41104 37612 41110 37664
rect 42886 37612 42892 37664
rect 42944 37652 42950 37664
rect 47394 37652 47400 37664
rect 42944 37624 47400 37652
rect 42944 37612 42950 37624
rect 47394 37612 47400 37624
rect 47452 37612 47458 37664
rect 47854 37652 47860 37664
rect 47815 37624 47860 37652
rect 47854 37612 47860 37624
rect 47912 37612 47918 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 24029 37451 24087 37457
rect 24029 37417 24041 37451
rect 24075 37448 24087 37451
rect 24762 37448 24768 37460
rect 24075 37420 24768 37448
rect 24075 37417 24087 37420
rect 24029 37411 24087 37417
rect 24762 37408 24768 37420
rect 24820 37408 24826 37460
rect 31018 37408 31024 37460
rect 31076 37448 31082 37460
rect 31665 37451 31723 37457
rect 31665 37448 31677 37451
rect 31076 37420 31677 37448
rect 31076 37408 31082 37420
rect 31665 37417 31677 37420
rect 31711 37448 31723 37451
rect 31711 37420 33088 37448
rect 31711 37417 31723 37420
rect 31665 37411 31723 37417
rect 33060 37392 33088 37420
rect 35434 37408 35440 37460
rect 35492 37448 35498 37460
rect 36173 37451 36231 37457
rect 35492 37420 35747 37448
rect 35492 37408 35498 37420
rect 25314 37380 25320 37392
rect 23676 37352 25320 37380
rect 23676 37321 23704 37352
rect 25314 37340 25320 37352
rect 25372 37380 25378 37392
rect 26050 37380 26056 37392
rect 25372 37352 26056 37380
rect 25372 37340 25378 37352
rect 26050 37340 26056 37352
rect 26108 37340 26114 37392
rect 26234 37380 26240 37392
rect 26195 37352 26240 37380
rect 26234 37340 26240 37352
rect 26292 37340 26298 37392
rect 33042 37380 33048 37392
rect 32955 37352 33048 37380
rect 33042 37340 33048 37352
rect 33100 37340 33106 37392
rect 34606 37340 34612 37392
rect 34664 37380 34670 37392
rect 34664 37352 35572 37380
rect 34664 37340 34670 37352
rect 35544 37324 35572 37352
rect 23661 37315 23719 37321
rect 23661 37281 23673 37315
rect 23707 37281 23719 37315
rect 23661 37275 23719 37281
rect 24581 37315 24639 37321
rect 24581 37281 24593 37315
rect 24627 37312 24639 37315
rect 24946 37312 24952 37324
rect 24627 37284 24952 37312
rect 24627 37281 24639 37284
rect 24581 37275 24639 37281
rect 24946 37272 24952 37284
rect 25004 37272 25010 37324
rect 26145 37315 26203 37321
rect 26145 37281 26157 37315
rect 26191 37312 26203 37315
rect 27522 37312 27528 37324
rect 26191 37284 27528 37312
rect 26191 37281 26203 37284
rect 26145 37275 26203 37281
rect 27522 37272 27528 37284
rect 27580 37272 27586 37324
rect 27982 37312 27988 37324
rect 27943 37284 27988 37312
rect 27982 37272 27988 37284
rect 28040 37272 28046 37324
rect 33597 37315 33655 37321
rect 33597 37281 33609 37315
rect 33643 37312 33655 37315
rect 34698 37312 34704 37324
rect 33643 37284 34704 37312
rect 33643 37281 33655 37284
rect 33597 37275 33655 37281
rect 34698 37272 34704 37284
rect 34756 37272 34762 37324
rect 35526 37312 35532 37324
rect 35487 37284 35532 37312
rect 35526 37272 35532 37284
rect 35584 37272 35590 37324
rect 23845 37247 23903 37253
rect 23845 37213 23857 37247
rect 23891 37244 23903 37247
rect 24670 37244 24676 37256
rect 23891 37216 24676 37244
rect 23891 37213 23903 37216
rect 23845 37207 23903 37213
rect 24670 37204 24676 37216
rect 24728 37244 24734 37256
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 24728 37216 24777 37244
rect 24728 37204 24734 37216
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 26050 37244 26056 37256
rect 26011 37216 26056 37244
rect 24765 37207 24823 37213
rect 26050 37204 26056 37216
rect 26108 37204 26114 37256
rect 26326 37244 26332 37256
rect 26287 37216 26332 37244
rect 26326 37204 26332 37216
rect 26384 37204 26390 37256
rect 28166 37244 28172 37256
rect 28127 37216 28172 37244
rect 28166 37204 28172 37216
rect 28224 37204 28230 37256
rect 30285 37247 30343 37253
rect 30285 37213 30297 37247
rect 30331 37244 30343 37247
rect 32122 37244 32128 37256
rect 30331 37216 32128 37244
rect 30331 37213 30343 37216
rect 30285 37207 30343 37213
rect 32122 37204 32128 37216
rect 32180 37204 32186 37256
rect 32306 37244 32312 37256
rect 32267 37216 32312 37244
rect 32306 37204 32312 37216
rect 32364 37204 32370 37256
rect 33318 37244 33324 37256
rect 33231 37216 33324 37244
rect 33318 37204 33324 37216
rect 33376 37244 33382 37256
rect 33962 37244 33968 37256
rect 33376 37216 33968 37244
rect 33376 37204 33382 37216
rect 33962 37204 33968 37216
rect 34020 37204 34026 37256
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35719 37244 35747 37420
rect 36173 37417 36185 37451
rect 36219 37448 36231 37451
rect 37274 37448 37280 37460
rect 36219 37420 37280 37448
rect 36219 37417 36231 37420
rect 36173 37411 36231 37417
rect 37274 37408 37280 37420
rect 37332 37408 37338 37460
rect 37918 37448 37924 37460
rect 37879 37420 37924 37448
rect 37918 37408 37924 37420
rect 37976 37448 37982 37460
rect 42794 37448 42800 37460
rect 37976 37420 42800 37448
rect 37976 37408 37982 37420
rect 42794 37408 42800 37420
rect 42852 37408 42858 37460
rect 45649 37451 45707 37457
rect 45649 37417 45661 37451
rect 45695 37417 45707 37451
rect 45649 37411 45707 37417
rect 45833 37451 45891 37457
rect 45833 37417 45845 37451
rect 45879 37448 45891 37451
rect 46290 37448 46296 37460
rect 45879 37420 46296 37448
rect 45879 37417 45891 37420
rect 45833 37411 45891 37417
rect 43441 37383 43499 37389
rect 43441 37349 43453 37383
rect 43487 37349 43499 37383
rect 45664 37380 45692 37411
rect 46290 37408 46296 37420
rect 46348 37408 46354 37460
rect 46198 37380 46204 37392
rect 45664 37352 46204 37380
rect 43441 37343 43499 37349
rect 40405 37315 40463 37321
rect 40405 37281 40417 37315
rect 40451 37312 40463 37315
rect 41046 37312 41052 37324
rect 40451 37284 41052 37312
rect 40451 37281 40463 37284
rect 40405 37275 40463 37281
rect 41046 37272 41052 37284
rect 41104 37272 41110 37324
rect 43456 37312 43484 37343
rect 46198 37340 46204 37352
rect 46256 37340 46262 37392
rect 43901 37315 43959 37321
rect 43901 37312 43913 37315
rect 43456 37284 43913 37312
rect 43901 37281 43913 37284
rect 43947 37312 43959 37315
rect 44174 37312 44180 37324
rect 43947 37284 44180 37312
rect 43947 37281 43959 37284
rect 43901 37275 43959 37281
rect 44174 37272 44180 37284
rect 44232 37272 44238 37324
rect 48222 37312 48228 37324
rect 48183 37284 48228 37312
rect 48222 37272 48228 37284
rect 48280 37272 48286 37324
rect 35989 37247 36047 37253
rect 35989 37244 36001 37247
rect 35719 37216 36001 37244
rect 35069 37207 35127 37213
rect 35989 37213 36001 37216
rect 36035 37213 36047 37247
rect 35989 37207 36047 37213
rect 36081 37247 36139 37253
rect 36081 37213 36093 37247
rect 36127 37244 36139 37247
rect 36814 37244 36820 37256
rect 36127 37216 36820 37244
rect 36127 37213 36139 37216
rect 36081 37207 36139 37213
rect 36814 37204 36820 37216
rect 36872 37204 36878 37256
rect 37182 37204 37188 37256
rect 37240 37244 37246 37256
rect 40034 37244 40040 37256
rect 37240 37216 40040 37244
rect 37240 37204 37246 37216
rect 40034 37204 40040 37216
rect 40092 37204 40098 37256
rect 40310 37244 40316 37256
rect 40271 37216 40316 37244
rect 40310 37204 40316 37216
rect 40368 37204 40374 37256
rect 41141 37247 41199 37253
rect 41141 37213 41153 37247
rect 41187 37213 41199 37247
rect 41141 37207 41199 37213
rect 42061 37247 42119 37253
rect 42061 37213 42073 37247
rect 42107 37244 42119 37247
rect 43346 37244 43352 37256
rect 42107 37216 43352 37244
rect 42107 37213 42119 37216
rect 42061 37207 42119 37213
rect 26602 37136 26608 37188
rect 26660 37176 26666 37188
rect 28902 37176 28908 37188
rect 26660 37148 28908 37176
rect 26660 37136 26666 37148
rect 28902 37136 28908 37148
rect 28960 37136 28966 37188
rect 30552 37179 30610 37185
rect 30552 37145 30564 37179
rect 30598 37176 30610 37179
rect 30598 37148 31754 37176
rect 30598 37145 30610 37148
rect 30552 37139 30610 37145
rect 23382 37068 23388 37120
rect 23440 37108 23446 37120
rect 24949 37111 25007 37117
rect 24949 37108 24961 37111
rect 23440 37080 24961 37108
rect 23440 37068 23446 37080
rect 24949 37077 24961 37080
rect 24995 37077 25007 37111
rect 24949 37071 25007 37077
rect 25869 37111 25927 37117
rect 25869 37077 25881 37111
rect 25915 37108 25927 37111
rect 26234 37108 26240 37120
rect 25915 37080 26240 37108
rect 25915 37077 25927 37080
rect 25869 37071 25927 37077
rect 26234 37068 26240 37080
rect 26292 37068 26298 37120
rect 28353 37111 28411 37117
rect 28353 37077 28365 37111
rect 28399 37108 28411 37111
rect 28442 37108 28448 37120
rect 28399 37080 28448 37108
rect 28399 37077 28411 37080
rect 28353 37071 28411 37077
rect 28442 37068 28448 37080
rect 28500 37068 28506 37120
rect 31726 37108 31754 37148
rect 33134 37136 33140 37188
rect 33192 37176 33198 37188
rect 33410 37176 33416 37188
rect 33192 37148 33416 37176
rect 33192 37136 33198 37148
rect 33410 37136 33416 37148
rect 33468 37136 33474 37188
rect 35161 37179 35219 37185
rect 35161 37145 35173 37179
rect 35207 37145 35219 37179
rect 35161 37139 35219 37145
rect 32125 37111 32183 37117
rect 32125 37108 32137 37111
rect 31726 37080 32137 37108
rect 32125 37077 32137 37080
rect 32171 37077 32183 37111
rect 33226 37108 33232 37120
rect 33187 37080 33232 37108
rect 32125 37071 32183 37077
rect 33226 37068 33232 37080
rect 33284 37068 33290 37120
rect 34882 37108 34888 37120
rect 34843 37080 34888 37108
rect 34882 37068 34888 37080
rect 34940 37068 34946 37120
rect 35176 37108 35204 37139
rect 35250 37136 35256 37188
rect 35308 37176 35314 37188
rect 35391 37179 35449 37185
rect 35308 37148 35353 37176
rect 35308 37136 35314 37148
rect 35391 37145 35403 37179
rect 35437 37176 35449 37179
rect 36170 37176 36176 37188
rect 35437 37148 36176 37176
rect 35437 37145 35449 37148
rect 35391 37139 35449 37145
rect 36170 37136 36176 37148
rect 36228 37136 36234 37188
rect 37550 37136 37556 37188
rect 37608 37176 37614 37188
rect 37829 37179 37887 37185
rect 37829 37176 37841 37179
rect 37608 37148 37841 37176
rect 37608 37136 37614 37148
rect 37829 37145 37841 37148
rect 37875 37145 37887 37179
rect 37829 37139 37887 37145
rect 39942 37136 39948 37188
rect 40000 37176 40006 37188
rect 40522 37179 40580 37185
rect 40522 37176 40534 37179
rect 40000 37148 40534 37176
rect 40000 37136 40006 37148
rect 40522 37145 40534 37148
rect 40568 37145 40580 37179
rect 40522 37139 40580 37145
rect 35894 37108 35900 37120
rect 35176 37080 35900 37108
rect 35894 37068 35900 37080
rect 35952 37068 35958 37120
rect 36357 37111 36415 37117
rect 36357 37077 36369 37111
rect 36403 37108 36415 37111
rect 36446 37108 36452 37120
rect 36403 37080 36452 37108
rect 36403 37077 36415 37080
rect 36357 37071 36415 37077
rect 36446 37068 36452 37080
rect 36504 37068 36510 37120
rect 40681 37111 40739 37117
rect 40681 37077 40693 37111
rect 40727 37108 40739 37111
rect 40954 37108 40960 37120
rect 40727 37080 40960 37108
rect 40727 37077 40739 37080
rect 40681 37071 40739 37077
rect 40954 37068 40960 37080
rect 41012 37068 41018 37120
rect 41156 37108 41184 37207
rect 43346 37204 43352 37216
rect 43404 37204 43410 37256
rect 44082 37244 44088 37256
rect 43995 37216 44088 37244
rect 44082 37204 44088 37216
rect 44140 37204 44146 37256
rect 44266 37244 44272 37256
rect 44227 37216 44272 37244
rect 44266 37204 44272 37216
rect 44324 37204 44330 37256
rect 46477 37247 46535 37253
rect 46477 37213 46489 37247
rect 46523 37213 46535 37247
rect 46477 37207 46535 37213
rect 41414 37136 41420 37188
rect 41472 37176 41478 37188
rect 42328 37179 42386 37185
rect 41472 37148 41517 37176
rect 41472 37136 41478 37148
rect 42328 37145 42340 37179
rect 42374 37176 42386 37179
rect 42610 37176 42616 37188
rect 42374 37148 42616 37176
rect 42374 37145 42386 37148
rect 42328 37139 42386 37145
rect 42610 37136 42616 37148
rect 42668 37136 42674 37188
rect 44100 37176 44128 37204
rect 45370 37176 45376 37188
rect 44100 37148 45376 37176
rect 44100 37108 44128 37148
rect 45370 37136 45376 37148
rect 45428 37176 45434 37188
rect 45465 37179 45523 37185
rect 45465 37176 45477 37179
rect 45428 37148 45477 37176
rect 45428 37136 45434 37148
rect 45465 37145 45477 37148
rect 45511 37145 45523 37179
rect 45465 37139 45523 37145
rect 41156 37080 44128 37108
rect 45675 37111 45733 37117
rect 45675 37077 45687 37111
rect 45721 37108 45733 37111
rect 45830 37108 45836 37120
rect 45721 37080 45836 37108
rect 45721 37077 45733 37080
rect 45675 37071 45733 37077
rect 45830 37068 45836 37080
rect 45888 37068 45894 37120
rect 46492 37108 46520 37207
rect 46661 37179 46719 37185
rect 46661 37145 46673 37179
rect 46707 37176 46719 37179
rect 47854 37176 47860 37188
rect 46707 37148 47860 37176
rect 46707 37145 46719 37148
rect 46661 37139 46719 37145
rect 47854 37136 47860 37148
rect 47912 37136 47918 37188
rect 47946 37108 47952 37120
rect 46492 37080 47952 37108
rect 47946 37068 47952 37080
rect 48004 37068 48010 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 25159 36907 25217 36913
rect 25159 36873 25171 36907
rect 25205 36904 25217 36907
rect 25958 36904 25964 36916
rect 25205 36876 25964 36904
rect 25205 36873 25217 36876
rect 25159 36867 25217 36873
rect 25958 36864 25964 36876
rect 26016 36864 26022 36916
rect 28166 36864 28172 36916
rect 28224 36904 28230 36916
rect 30469 36907 30527 36913
rect 30469 36904 30481 36907
rect 28224 36876 30481 36904
rect 28224 36864 28230 36876
rect 30469 36873 30481 36876
rect 30515 36873 30527 36907
rect 30469 36867 30527 36873
rect 31757 36907 31815 36913
rect 31757 36873 31769 36907
rect 31803 36904 31815 36907
rect 32306 36904 32312 36916
rect 31803 36876 32312 36904
rect 31803 36873 31815 36876
rect 31757 36867 31815 36873
rect 24946 36836 24952 36848
rect 24859 36808 24952 36836
rect 24946 36796 24952 36808
rect 25004 36836 25010 36848
rect 25774 36836 25780 36848
rect 25004 36808 25780 36836
rect 25004 36796 25010 36808
rect 25774 36796 25780 36808
rect 25832 36796 25838 36848
rect 26142 36836 26148 36848
rect 26103 36808 26148 36836
rect 26142 36796 26148 36808
rect 26200 36796 26206 36848
rect 26234 36796 26240 36848
rect 26292 36845 26298 36848
rect 26292 36839 26321 36845
rect 26309 36805 26321 36839
rect 26292 36799 26321 36805
rect 26292 36796 26298 36799
rect 26970 36796 26976 36848
rect 27028 36836 27034 36848
rect 30484 36836 30512 36867
rect 32306 36864 32312 36876
rect 32364 36864 32370 36916
rect 35713 36907 35771 36913
rect 35713 36873 35725 36907
rect 35759 36873 35771 36907
rect 36170 36904 36176 36916
rect 36131 36876 36176 36904
rect 35713 36867 35771 36873
rect 32030 36836 32036 36848
rect 27028 36808 29132 36836
rect 30484 36808 32036 36836
rect 27028 36796 27034 36808
rect 24305 36771 24363 36777
rect 24305 36737 24317 36771
rect 24351 36768 24363 36771
rect 24670 36768 24676 36780
rect 24351 36740 24676 36768
rect 24351 36737 24363 36740
rect 24305 36731 24363 36737
rect 24670 36728 24676 36740
rect 24728 36728 24734 36780
rect 25961 36771 26019 36777
rect 25961 36768 25973 36771
rect 25332 36740 25973 36768
rect 24121 36703 24179 36709
rect 24121 36669 24133 36703
rect 24167 36700 24179 36703
rect 24167 36672 25176 36700
rect 24167 36669 24179 36672
rect 24121 36663 24179 36669
rect 24026 36524 24032 36576
rect 24084 36564 24090 36576
rect 25148 36573 25176 36672
rect 25332 36641 25360 36740
rect 25961 36737 25973 36740
rect 26007 36737 26019 36771
rect 25961 36731 26019 36737
rect 26053 36771 26111 36777
rect 26053 36737 26065 36771
rect 26099 36737 26111 36771
rect 27424 36771 27482 36777
rect 27424 36768 27436 36771
rect 26053 36731 26111 36737
rect 26206 36740 27436 36768
rect 26068 36700 26096 36731
rect 26206 36700 26234 36740
rect 27424 36737 27436 36740
rect 27470 36768 27482 36771
rect 28258 36768 28264 36780
rect 27470 36740 28264 36768
rect 27470 36737 27482 36740
rect 27424 36731 27482 36737
rect 28258 36728 28264 36740
rect 28316 36728 28322 36780
rect 26068 36672 26234 36700
rect 26421 36703 26479 36709
rect 26421 36669 26433 36703
rect 26467 36700 26479 36703
rect 26602 36700 26608 36712
rect 26467 36672 26608 36700
rect 26467 36669 26479 36672
rect 26421 36663 26479 36669
rect 26602 36660 26608 36672
rect 26660 36660 26666 36712
rect 27154 36700 27160 36712
rect 27115 36672 27160 36700
rect 27154 36660 27160 36672
rect 27212 36660 27218 36712
rect 25317 36635 25375 36641
rect 25317 36601 25329 36635
rect 25363 36601 25375 36635
rect 26050 36632 26056 36644
rect 25317 36595 25375 36601
rect 25424 36604 26056 36632
rect 24489 36567 24547 36573
rect 24489 36564 24501 36567
rect 24084 36536 24501 36564
rect 24084 36524 24090 36536
rect 24489 36533 24501 36536
rect 24535 36533 24547 36567
rect 24489 36527 24547 36533
rect 25133 36567 25191 36573
rect 25133 36533 25145 36567
rect 25179 36564 25191 36567
rect 25424 36564 25452 36604
rect 26050 36592 26056 36604
rect 26108 36592 26114 36644
rect 25774 36564 25780 36576
rect 25179 36536 25452 36564
rect 25735 36536 25780 36564
rect 25179 36533 25191 36536
rect 25133 36527 25191 36533
rect 25774 36524 25780 36536
rect 25832 36524 25838 36576
rect 25866 36524 25872 36576
rect 25924 36564 25930 36576
rect 27338 36564 27344 36576
rect 25924 36536 27344 36564
rect 25924 36524 25930 36536
rect 27338 36524 27344 36536
rect 27396 36564 27402 36576
rect 28537 36567 28595 36573
rect 28537 36564 28549 36567
rect 27396 36536 28549 36564
rect 27396 36524 27402 36536
rect 28537 36533 28549 36536
rect 28583 36533 28595 36567
rect 29104 36564 29132 36808
rect 32030 36796 32036 36808
rect 32088 36796 32094 36848
rect 32122 36796 32128 36848
rect 32180 36836 32186 36848
rect 34600 36839 34658 36845
rect 32180 36808 34376 36836
rect 32180 36796 32186 36808
rect 30377 36771 30435 36777
rect 30377 36737 30389 36771
rect 30423 36768 30435 36771
rect 30650 36768 30656 36780
rect 30423 36740 30656 36768
rect 30423 36737 30435 36740
rect 30377 36731 30435 36737
rect 30650 36728 30656 36740
rect 30708 36728 30714 36780
rect 31202 36728 31208 36780
rect 31260 36768 31266 36780
rect 31573 36771 31631 36777
rect 31573 36768 31585 36771
rect 31260 36740 31585 36768
rect 31260 36728 31266 36740
rect 31573 36737 31585 36740
rect 31619 36737 31631 36771
rect 33134 36768 33140 36780
rect 33095 36740 33140 36768
rect 31573 36731 31631 36737
rect 33134 36728 33140 36740
rect 33192 36728 33198 36780
rect 33318 36768 33324 36780
rect 33279 36740 33324 36768
rect 33318 36728 33324 36740
rect 33376 36728 33382 36780
rect 34348 36777 34376 36808
rect 34600 36805 34612 36839
rect 34646 36836 34658 36839
rect 34882 36836 34888 36848
rect 34646 36808 34888 36836
rect 34646 36805 34658 36808
rect 34600 36799 34658 36805
rect 34882 36796 34888 36808
rect 34940 36796 34946 36848
rect 35618 36796 35624 36848
rect 35676 36836 35682 36848
rect 35728 36836 35756 36867
rect 36170 36864 36176 36876
rect 36228 36864 36234 36916
rect 37458 36864 37464 36916
rect 37516 36904 37522 36916
rect 40313 36907 40371 36913
rect 40313 36904 40325 36907
rect 37516 36876 40325 36904
rect 37516 36864 37522 36876
rect 40313 36873 40325 36876
rect 40359 36873 40371 36907
rect 42610 36904 42616 36916
rect 42571 36876 42616 36904
rect 40313 36867 40371 36873
rect 42610 36864 42616 36876
rect 42668 36864 42674 36916
rect 35676 36808 36676 36836
rect 35676 36796 35682 36808
rect 33413 36771 33471 36777
rect 33413 36737 33425 36771
rect 33459 36737 33471 36771
rect 33413 36731 33471 36737
rect 34333 36771 34391 36777
rect 34333 36737 34345 36771
rect 34379 36737 34391 36771
rect 34333 36731 34391 36737
rect 31389 36703 31447 36709
rect 31389 36669 31401 36703
rect 31435 36700 31447 36703
rect 31435 36672 31754 36700
rect 31435 36669 31447 36672
rect 31389 36663 31447 36669
rect 31726 36632 31754 36672
rect 33042 36660 33048 36712
rect 33100 36700 33106 36712
rect 33428 36700 33456 36731
rect 35342 36728 35348 36780
rect 35400 36768 35406 36780
rect 36357 36771 36415 36777
rect 36357 36768 36369 36771
rect 35400 36740 36369 36768
rect 35400 36728 35406 36740
rect 36357 36737 36369 36740
rect 36403 36737 36415 36771
rect 36357 36731 36415 36737
rect 36446 36728 36452 36780
rect 36504 36768 36510 36780
rect 36648 36777 36676 36808
rect 36722 36796 36728 36848
rect 36780 36836 36786 36848
rect 39022 36836 39028 36848
rect 36780 36808 39028 36836
rect 36780 36796 36786 36808
rect 39022 36796 39028 36808
rect 39080 36796 39086 36848
rect 39206 36796 39212 36848
rect 39264 36836 39270 36848
rect 47670 36836 47676 36848
rect 39264 36808 47676 36836
rect 39264 36796 39270 36808
rect 47670 36796 47676 36808
rect 47728 36836 47734 36848
rect 47728 36808 47808 36836
rect 47728 36796 47734 36808
rect 36633 36771 36691 36777
rect 36504 36740 36549 36768
rect 36504 36728 36510 36740
rect 36633 36737 36645 36771
rect 36679 36737 36691 36771
rect 36633 36731 36691 36737
rect 37550 36728 37556 36780
rect 37608 36768 37614 36780
rect 37645 36771 37703 36777
rect 37645 36768 37657 36771
rect 37608 36740 37657 36768
rect 37608 36728 37614 36740
rect 37645 36737 37657 36740
rect 37691 36737 37703 36771
rect 37645 36731 37703 36737
rect 41046 36728 41052 36780
rect 41104 36768 41110 36780
rect 41417 36771 41475 36777
rect 41417 36768 41429 36771
rect 41104 36740 41429 36768
rect 41104 36728 41110 36740
rect 41417 36737 41429 36740
rect 41463 36737 41475 36771
rect 42794 36768 42800 36780
rect 42755 36740 42800 36768
rect 41417 36731 41475 36737
rect 42794 36728 42800 36740
rect 42852 36728 42858 36780
rect 47780 36777 47808 36808
rect 47765 36771 47823 36777
rect 47765 36737 47777 36771
rect 47811 36737 47823 36771
rect 47765 36731 47823 36737
rect 33100 36672 33456 36700
rect 33100 36660 33106 36672
rect 37274 36660 37280 36712
rect 37332 36700 37338 36712
rect 37461 36703 37519 36709
rect 37461 36700 37473 36703
rect 37332 36672 37473 36700
rect 37332 36660 37338 36672
rect 37461 36669 37473 36672
rect 37507 36700 37519 36703
rect 38562 36700 38568 36712
rect 37507 36672 38568 36700
rect 37507 36669 37519 36672
rect 37461 36663 37519 36669
rect 38562 36660 38568 36672
rect 38620 36660 38626 36712
rect 40310 36660 40316 36712
rect 40368 36700 40374 36712
rect 41138 36700 41144 36712
rect 40368 36672 41144 36700
rect 40368 36660 40374 36672
rect 41138 36660 41144 36672
rect 41196 36700 41202 36712
rect 41233 36703 41291 36709
rect 41233 36700 41245 36703
rect 41196 36672 41245 36700
rect 41196 36660 41202 36672
rect 41233 36669 41245 36672
rect 41279 36669 41291 36703
rect 41233 36663 41291 36669
rect 36541 36635 36599 36641
rect 36541 36632 36553 36635
rect 31726 36604 33272 36632
rect 33244 36576 33272 36604
rect 35268 36604 36553 36632
rect 33134 36564 33140 36576
rect 29104 36536 33140 36564
rect 28537 36527 28595 36533
rect 33134 36524 33140 36536
rect 33192 36524 33198 36576
rect 33226 36524 33232 36576
rect 33284 36564 33290 36576
rect 33410 36564 33416 36576
rect 33284 36536 33416 36564
rect 33284 36524 33290 36536
rect 33410 36524 33416 36536
rect 33468 36524 33474 36576
rect 33597 36567 33655 36573
rect 33597 36533 33609 36567
rect 33643 36564 33655 36567
rect 35268 36564 35296 36604
rect 36541 36601 36553 36604
rect 36587 36601 36599 36635
rect 36541 36595 36599 36601
rect 37826 36564 37832 36576
rect 33643 36536 35296 36564
rect 37787 36536 37832 36564
rect 33643 36533 33655 36536
rect 33597 36527 33655 36533
rect 37826 36524 37832 36536
rect 37884 36524 37890 36576
rect 39666 36524 39672 36576
rect 39724 36564 39730 36576
rect 41601 36567 41659 36573
rect 41601 36564 41613 36567
rect 39724 36536 41613 36564
rect 39724 36524 39730 36536
rect 41601 36533 41613 36536
rect 41647 36533 41659 36567
rect 41601 36527 41659 36533
rect 46474 36524 46480 36576
rect 46532 36564 46538 36576
rect 47213 36567 47271 36573
rect 47213 36564 47225 36567
rect 46532 36536 47225 36564
rect 46532 36524 46538 36536
rect 47213 36533 47225 36536
rect 47259 36533 47271 36567
rect 47854 36564 47860 36576
rect 47815 36536 47860 36564
rect 47213 36527 47271 36533
rect 47854 36524 47860 36536
rect 47912 36524 47918 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 28258 36360 28264 36372
rect 28219 36332 28264 36360
rect 28258 36320 28264 36332
rect 28316 36320 28322 36372
rect 32122 36320 32128 36372
rect 32180 36360 32186 36372
rect 32493 36363 32551 36369
rect 32493 36360 32505 36363
rect 32180 36332 32505 36360
rect 32180 36320 32186 36332
rect 32493 36329 32505 36332
rect 32539 36329 32551 36363
rect 32493 36323 32551 36329
rect 33134 36320 33140 36372
rect 33192 36360 33198 36372
rect 39206 36360 39212 36372
rect 33192 36332 39212 36360
rect 33192 36320 33198 36332
rect 39206 36320 39212 36332
rect 39264 36320 39270 36372
rect 39117 36295 39175 36301
rect 39117 36261 39129 36295
rect 39163 36292 39175 36295
rect 39942 36292 39948 36304
rect 39163 36264 39948 36292
rect 39163 36261 39175 36264
rect 39117 36255 39175 36261
rect 39942 36252 39948 36264
rect 40000 36252 40006 36304
rect 40034 36252 40040 36304
rect 40092 36292 40098 36304
rect 40313 36295 40371 36301
rect 40313 36292 40325 36295
rect 40092 36264 40325 36292
rect 40092 36252 40098 36264
rect 40313 36261 40325 36264
rect 40359 36261 40371 36295
rect 40313 36255 40371 36261
rect 37182 36184 37188 36236
rect 37240 36224 37246 36236
rect 38841 36227 38899 36233
rect 38841 36224 38853 36227
rect 37240 36196 38853 36224
rect 37240 36184 37246 36196
rect 38841 36193 38853 36196
rect 38887 36193 38899 36227
rect 38841 36187 38899 36193
rect 39022 36184 39028 36236
rect 39080 36224 39086 36236
rect 46474 36224 46480 36236
rect 39080 36196 41414 36224
rect 46435 36196 46480 36224
rect 39080 36184 39086 36196
rect 23382 36156 23388 36168
rect 23343 36128 23388 36156
rect 23382 36116 23388 36128
rect 23440 36116 23446 36168
rect 24026 36156 24032 36168
rect 23987 36128 24032 36156
rect 24026 36116 24032 36128
rect 24084 36116 24090 36168
rect 28442 36156 28448 36168
rect 28403 36128 28448 36156
rect 28442 36116 28448 36128
rect 28500 36116 28506 36168
rect 34514 36116 34520 36168
rect 34572 36156 34578 36168
rect 35437 36159 35495 36165
rect 35437 36156 35449 36159
rect 34572 36128 35449 36156
rect 34572 36116 34578 36128
rect 35437 36125 35449 36128
rect 35483 36156 35495 36159
rect 37458 36156 37464 36168
rect 35483 36128 37464 36156
rect 35483 36125 35495 36128
rect 35437 36119 35495 36125
rect 37458 36116 37464 36128
rect 37516 36116 37522 36168
rect 39942 36116 39948 36168
rect 40000 36156 40006 36168
rect 40037 36159 40095 36165
rect 40037 36156 40049 36159
rect 40000 36128 40049 36156
rect 40000 36116 40006 36128
rect 40037 36125 40049 36128
rect 40083 36125 40095 36159
rect 40037 36119 40095 36125
rect 40957 36159 41015 36165
rect 40957 36125 40969 36159
rect 41003 36156 41015 36159
rect 41046 36156 41052 36168
rect 41003 36128 41052 36156
rect 41003 36125 41015 36128
rect 40957 36119 41015 36125
rect 41046 36116 41052 36128
rect 41104 36116 41110 36168
rect 41138 36116 41144 36168
rect 41196 36156 41202 36168
rect 41386 36156 41414 36196
rect 46474 36184 46480 36196
rect 46532 36184 46538 36236
rect 46661 36227 46719 36233
rect 46661 36193 46673 36227
rect 46707 36224 46719 36227
rect 47854 36224 47860 36236
rect 46707 36196 47860 36224
rect 46707 36193 46719 36196
rect 46661 36187 46719 36193
rect 47854 36184 47860 36196
rect 47912 36184 47918 36236
rect 48222 36224 48228 36236
rect 48183 36196 48228 36224
rect 48222 36184 48228 36196
rect 48280 36184 48286 36236
rect 41601 36159 41659 36165
rect 41601 36156 41613 36159
rect 41196 36128 41241 36156
rect 41386 36128 41613 36156
rect 41196 36116 41202 36128
rect 41601 36125 41613 36128
rect 41647 36125 41659 36159
rect 41601 36119 41659 36125
rect 44085 36159 44143 36165
rect 44085 36125 44097 36159
rect 44131 36156 44143 36159
rect 44174 36156 44180 36168
rect 44131 36128 44180 36156
rect 44131 36125 44143 36128
rect 44085 36119 44143 36125
rect 44174 36116 44180 36128
rect 44232 36116 44238 36168
rect 44269 36159 44327 36165
rect 44269 36125 44281 36159
rect 44315 36125 44327 36159
rect 44269 36119 44327 36125
rect 26053 36091 26111 36097
rect 26053 36057 26065 36091
rect 26099 36088 26111 36091
rect 31205 36091 31263 36097
rect 31205 36088 31217 36091
rect 26099 36060 31217 36088
rect 26099 36057 26111 36060
rect 26053 36051 26111 36057
rect 31205 36057 31217 36060
rect 31251 36088 31263 36091
rect 35704 36091 35762 36097
rect 31251 36060 31754 36088
rect 31251 36057 31263 36060
rect 31205 36051 31263 36057
rect 23201 36023 23259 36029
rect 23201 35989 23213 36023
rect 23247 36020 23259 36023
rect 23750 36020 23756 36032
rect 23247 35992 23756 36020
rect 23247 35989 23259 35992
rect 23201 35983 23259 35989
rect 23750 35980 23756 35992
rect 23808 35980 23814 36032
rect 23845 36023 23903 36029
rect 23845 35989 23857 36023
rect 23891 36020 23903 36023
rect 24026 36020 24032 36032
rect 23891 35992 24032 36020
rect 23891 35989 23903 35992
rect 23845 35983 23903 35989
rect 24026 35980 24032 35992
rect 24084 35980 24090 36032
rect 26234 35980 26240 36032
rect 26292 36020 26298 36032
rect 27154 36020 27160 36032
rect 26292 35992 27160 36020
rect 26292 35980 26298 35992
rect 27154 35980 27160 35992
rect 27212 36020 27218 36032
rect 27341 36023 27399 36029
rect 27341 36020 27353 36023
rect 27212 35992 27353 36020
rect 27212 35980 27218 35992
rect 27341 35989 27353 35992
rect 27387 35989 27399 36023
rect 31726 36020 31754 36060
rect 35704 36057 35716 36091
rect 35750 36088 35762 36091
rect 35894 36088 35900 36100
rect 35750 36060 35900 36088
rect 35750 36057 35762 36060
rect 35704 36051 35762 36057
rect 35894 36048 35900 36060
rect 35952 36048 35958 36100
rect 43346 36088 43352 36100
rect 43307 36060 43352 36088
rect 43346 36048 43352 36060
rect 43404 36048 43410 36100
rect 43990 36048 43996 36100
rect 44048 36088 44054 36100
rect 44284 36088 44312 36119
rect 44048 36060 44312 36088
rect 44048 36048 44054 36060
rect 36722 36020 36728 36032
rect 31726 35992 36728 36020
rect 27341 35983 27399 35989
rect 36722 35980 36728 35992
rect 36780 35980 36786 36032
rect 36814 35980 36820 36032
rect 36872 36020 36878 36032
rect 39301 36023 39359 36029
rect 36872 35992 36917 36020
rect 36872 35980 36878 35992
rect 39301 35989 39313 36023
rect 39347 36020 39359 36023
rect 39574 36020 39580 36032
rect 39347 35992 39580 36020
rect 39347 35989 39359 35992
rect 39301 35983 39359 35989
rect 39574 35980 39580 35992
rect 39632 35980 39638 36032
rect 40494 36020 40500 36032
rect 40455 35992 40500 36020
rect 40494 35980 40500 35992
rect 40552 35980 40558 36032
rect 40678 35980 40684 36032
rect 40736 36020 40742 36032
rect 41049 36023 41107 36029
rect 41049 36020 41061 36023
rect 40736 35992 41061 36020
rect 40736 35980 40742 35992
rect 41049 35989 41061 35992
rect 41095 35989 41107 36023
rect 44174 36020 44180 36032
rect 44135 35992 44180 36020
rect 41049 35983 41107 35989
rect 44174 35980 44180 35992
rect 44232 35980 44238 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 25958 35816 25964 35828
rect 25919 35788 25964 35816
rect 25958 35776 25964 35788
rect 26016 35776 26022 35828
rect 27522 35816 27528 35828
rect 27483 35788 27528 35816
rect 27522 35776 27528 35788
rect 27580 35776 27586 35828
rect 33410 35776 33416 35828
rect 33468 35816 33474 35828
rect 33689 35819 33747 35825
rect 33689 35816 33701 35819
rect 33468 35788 33701 35816
rect 33468 35776 33474 35788
rect 33689 35785 33701 35788
rect 33735 35785 33747 35819
rect 33689 35779 33747 35785
rect 34698 35776 34704 35828
rect 34756 35825 34762 35828
rect 34756 35819 34775 35825
rect 34763 35785 34775 35819
rect 34882 35816 34888 35828
rect 34843 35788 34888 35816
rect 34756 35779 34775 35785
rect 34756 35776 34762 35779
rect 34882 35776 34888 35788
rect 34940 35776 34946 35828
rect 35894 35816 35900 35828
rect 35855 35788 35900 35816
rect 35894 35776 35900 35788
rect 35952 35776 35958 35828
rect 39482 35816 39488 35828
rect 38764 35788 39488 35816
rect 23750 35708 23756 35760
rect 23808 35748 23814 35760
rect 24826 35751 24884 35757
rect 24826 35748 24838 35751
rect 23808 35720 24838 35748
rect 23808 35708 23814 35720
rect 24826 35717 24838 35720
rect 24872 35717 24884 35751
rect 24826 35711 24884 35717
rect 34517 35751 34575 35757
rect 34517 35717 34529 35751
rect 34563 35748 34575 35751
rect 36814 35748 36820 35760
rect 34563 35720 36820 35748
rect 34563 35717 34575 35720
rect 34517 35711 34575 35717
rect 25314 35640 25320 35692
rect 25372 35680 25378 35692
rect 27157 35683 27215 35689
rect 27157 35680 27169 35683
rect 25372 35652 27169 35680
rect 25372 35640 25378 35652
rect 27157 35649 27169 35652
rect 27203 35649 27215 35683
rect 27338 35680 27344 35692
rect 27299 35652 27344 35680
rect 27157 35643 27215 35649
rect 27338 35640 27344 35652
rect 27396 35640 27402 35692
rect 28074 35640 28080 35692
rect 28132 35680 28138 35692
rect 29181 35683 29239 35689
rect 29181 35680 29193 35683
rect 28132 35652 29193 35680
rect 28132 35640 28138 35652
rect 29181 35649 29193 35652
rect 29227 35649 29239 35683
rect 29181 35643 29239 35649
rect 29270 35640 29276 35692
rect 29328 35680 29334 35692
rect 29437 35683 29495 35689
rect 29437 35680 29449 35683
rect 29328 35652 29449 35680
rect 29328 35640 29334 35652
rect 29437 35649 29449 35652
rect 29483 35649 29495 35683
rect 29437 35643 29495 35649
rect 32122 35640 32128 35692
rect 32180 35680 32186 35692
rect 32582 35689 32588 35692
rect 32309 35683 32367 35689
rect 32309 35680 32321 35683
rect 32180 35652 32321 35680
rect 32180 35640 32186 35652
rect 32309 35649 32321 35652
rect 32355 35649 32367 35683
rect 32309 35643 32367 35649
rect 32576 35643 32588 35689
rect 32640 35680 32646 35692
rect 32640 35652 32676 35680
rect 32582 35640 32588 35643
rect 32640 35640 32646 35652
rect 33686 35640 33692 35692
rect 33744 35680 33750 35692
rect 34532 35680 34560 35711
rect 36814 35708 36820 35720
rect 36872 35708 36878 35760
rect 33744 35652 34560 35680
rect 36081 35683 36139 35689
rect 33744 35640 33750 35652
rect 36081 35649 36093 35683
rect 36127 35680 36139 35683
rect 37826 35680 37832 35692
rect 36127 35652 37832 35680
rect 36127 35649 36139 35652
rect 36081 35643 36139 35649
rect 37826 35640 37832 35652
rect 37884 35640 37890 35692
rect 38473 35683 38531 35689
rect 38473 35649 38485 35683
rect 38519 35649 38531 35683
rect 38473 35643 38531 35649
rect 38565 35683 38623 35689
rect 38565 35649 38577 35683
rect 38611 35680 38623 35683
rect 38764 35680 38792 35788
rect 39482 35776 39488 35788
rect 39540 35816 39546 35828
rect 40678 35816 40684 35828
rect 39540 35788 40684 35816
rect 39540 35776 39546 35788
rect 40678 35776 40684 35788
rect 40736 35776 40742 35828
rect 41322 35776 41328 35828
rect 41380 35816 41386 35828
rect 41877 35819 41935 35825
rect 41380 35776 41414 35816
rect 41877 35785 41889 35819
rect 41923 35816 41935 35819
rect 42794 35816 42800 35828
rect 41923 35788 42800 35816
rect 41923 35785 41935 35788
rect 41877 35779 41935 35785
rect 42794 35776 42800 35788
rect 42852 35776 42858 35828
rect 43254 35776 43260 35828
rect 43312 35816 43318 35828
rect 43312 35788 43484 35816
rect 43312 35776 43318 35788
rect 40494 35748 40500 35760
rect 38856 35720 40500 35748
rect 38856 35689 38884 35720
rect 38611 35652 38792 35680
rect 38841 35683 38899 35689
rect 38611 35649 38623 35652
rect 38565 35643 38623 35649
rect 38841 35649 38853 35683
rect 38887 35649 38899 35683
rect 39298 35680 39304 35692
rect 39259 35652 39304 35680
rect 38841 35643 38899 35649
rect 24578 35612 24584 35624
rect 24539 35584 24584 35612
rect 24578 35572 24584 35584
rect 24636 35572 24642 35624
rect 38488 35544 38516 35643
rect 39298 35640 39304 35652
rect 39356 35640 39362 35692
rect 39482 35680 39488 35692
rect 39443 35652 39488 35680
rect 39482 35640 39488 35652
rect 39540 35640 39546 35692
rect 39574 35640 39580 35692
rect 39632 35680 39638 35692
rect 39868 35689 39896 35720
rect 40494 35708 40500 35720
rect 40552 35748 40558 35760
rect 40552 35720 40816 35748
rect 40552 35708 40558 35720
rect 39853 35683 39911 35689
rect 39632 35652 39677 35680
rect 39632 35640 39638 35652
rect 39853 35649 39865 35683
rect 39899 35649 39911 35683
rect 40678 35680 40684 35692
rect 40639 35652 40684 35680
rect 39853 35643 39911 35649
rect 40678 35640 40684 35652
rect 40736 35640 40742 35692
rect 40788 35689 40816 35720
rect 40773 35683 40831 35689
rect 40773 35649 40785 35683
rect 40819 35649 40831 35683
rect 40954 35680 40960 35692
rect 40915 35652 40960 35680
rect 40773 35643 40831 35649
rect 40954 35640 40960 35652
rect 41012 35640 41018 35692
rect 41046 35640 41052 35692
rect 41104 35680 41110 35692
rect 41386 35680 41414 35776
rect 43346 35748 43352 35760
rect 42812 35720 43352 35748
rect 42812 35689 42840 35720
rect 43346 35708 43352 35720
rect 43404 35708 43410 35760
rect 43456 35748 43484 35788
rect 44266 35776 44272 35828
rect 44324 35816 44330 35828
rect 45005 35819 45063 35825
rect 45005 35816 45017 35819
rect 44324 35788 45017 35816
rect 44324 35776 44330 35788
rect 45005 35785 45017 35788
rect 45051 35785 45063 35819
rect 45005 35779 45063 35785
rect 46845 35751 46903 35757
rect 46845 35748 46857 35751
rect 43456 35720 46857 35748
rect 46845 35717 46857 35720
rect 46891 35748 46903 35751
rect 47118 35748 47124 35760
rect 46891 35720 47124 35748
rect 46891 35717 46903 35720
rect 46845 35711 46903 35717
rect 47118 35708 47124 35720
rect 47176 35708 47182 35760
rect 41509 35683 41567 35689
rect 41509 35680 41521 35683
rect 41104 35652 41149 35680
rect 41386 35652 41521 35680
rect 41104 35640 41110 35652
rect 41509 35649 41521 35652
rect 41555 35649 41567 35683
rect 41509 35643 41567 35649
rect 41693 35683 41751 35689
rect 41693 35649 41705 35683
rect 41739 35649 41751 35683
rect 41693 35643 41751 35649
rect 42797 35683 42855 35689
rect 42797 35649 42809 35683
rect 42843 35649 42855 35683
rect 42797 35643 42855 35649
rect 38749 35615 38807 35621
rect 38749 35581 38761 35615
rect 38795 35612 38807 35615
rect 39592 35612 39620 35640
rect 38795 35584 39620 35612
rect 38795 35581 38807 35584
rect 38749 35575 38807 35581
rect 39666 35572 39672 35624
rect 39724 35612 39730 35624
rect 39724 35584 39769 35612
rect 39724 35572 39730 35584
rect 39684 35544 39712 35572
rect 41046 35544 41052 35556
rect 38488 35516 39712 35544
rect 39776 35516 41052 35544
rect 27341 35479 27399 35485
rect 27341 35445 27353 35479
rect 27387 35476 27399 35479
rect 27982 35476 27988 35488
rect 27387 35448 27988 35476
rect 27387 35445 27399 35448
rect 27341 35439 27399 35445
rect 27982 35436 27988 35448
rect 28040 35436 28046 35488
rect 30558 35476 30564 35488
rect 30519 35448 30564 35476
rect 30558 35436 30564 35448
rect 30616 35436 30622 35488
rect 34701 35479 34759 35485
rect 34701 35445 34713 35479
rect 34747 35476 34759 35479
rect 34790 35476 34796 35488
rect 34747 35448 34796 35476
rect 34747 35445 34759 35448
rect 34701 35439 34759 35445
rect 34790 35436 34796 35448
rect 34848 35476 34854 35488
rect 35342 35476 35348 35488
rect 34848 35448 35348 35476
rect 34848 35436 34854 35448
rect 35342 35436 35348 35448
rect 35400 35436 35406 35488
rect 38289 35479 38347 35485
rect 38289 35445 38301 35479
rect 38335 35476 38347 35479
rect 38562 35476 38568 35488
rect 38335 35448 38568 35476
rect 38335 35445 38347 35448
rect 38289 35439 38347 35445
rect 38562 35436 38568 35448
rect 38620 35436 38626 35488
rect 39298 35436 39304 35488
rect 39356 35476 39362 35488
rect 39776 35476 39804 35516
rect 41046 35504 41052 35516
rect 41104 35504 41110 35556
rect 40034 35476 40040 35488
rect 39356 35448 39804 35476
rect 39995 35448 40040 35476
rect 39356 35436 39362 35448
rect 40034 35436 40040 35448
rect 40092 35436 40098 35488
rect 40494 35476 40500 35488
rect 40455 35448 40500 35476
rect 40494 35436 40500 35448
rect 40552 35436 40558 35488
rect 41708 35476 41736 35643
rect 42886 35640 42892 35692
rect 42944 35680 42950 35692
rect 43053 35683 43111 35689
rect 43053 35680 43065 35683
rect 42944 35652 43065 35680
rect 42944 35640 42950 35652
rect 43053 35649 43065 35652
rect 43099 35649 43111 35683
rect 43053 35643 43111 35649
rect 44821 35683 44879 35689
rect 44821 35649 44833 35683
rect 44867 35680 44879 35683
rect 45186 35680 45192 35692
rect 44867 35652 45192 35680
rect 44867 35649 44879 35652
rect 44821 35643 44879 35649
rect 45186 35640 45192 35652
rect 45244 35640 45250 35692
rect 46658 35680 46664 35692
rect 46619 35652 46664 35680
rect 46658 35640 46664 35652
rect 46716 35640 46722 35692
rect 46937 35683 46995 35689
rect 46937 35649 46949 35683
rect 46983 35680 46995 35683
rect 47210 35680 47216 35692
rect 46983 35652 47216 35680
rect 46983 35649 46995 35652
rect 46937 35643 46995 35649
rect 47210 35640 47216 35652
rect 47268 35640 47274 35692
rect 44358 35572 44364 35624
rect 44416 35612 44422 35624
rect 44637 35615 44695 35621
rect 44637 35612 44649 35615
rect 44416 35584 44649 35612
rect 44416 35572 44422 35584
rect 44637 35581 44649 35584
rect 44683 35581 44695 35615
rect 44637 35575 44695 35581
rect 48130 35544 48136 35556
rect 44100 35516 48136 35544
rect 44100 35476 44128 35516
rect 48130 35504 48136 35516
rect 48188 35504 48194 35556
rect 41708 35448 44128 35476
rect 44177 35479 44235 35485
rect 44177 35445 44189 35479
rect 44223 35476 44235 35479
rect 44358 35476 44364 35488
rect 44223 35448 44364 35476
rect 44223 35445 44235 35448
rect 44177 35439 44235 35445
rect 44358 35436 44364 35448
rect 44416 35436 44422 35488
rect 46661 35479 46719 35485
rect 46661 35445 46673 35479
rect 46707 35476 46719 35479
rect 47026 35476 47032 35488
rect 46707 35448 47032 35476
rect 46707 35445 46719 35448
rect 46661 35439 46719 35445
rect 47026 35436 47032 35448
rect 47084 35436 47090 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 26326 35232 26332 35284
rect 26384 35272 26390 35284
rect 26694 35272 26700 35284
rect 26384 35244 26700 35272
rect 26384 35232 26390 35244
rect 26694 35232 26700 35244
rect 26752 35272 26758 35284
rect 26973 35275 27031 35281
rect 26973 35272 26985 35275
rect 26752 35244 26985 35272
rect 26752 35232 26758 35244
rect 26973 35241 26985 35244
rect 27019 35241 27031 35275
rect 26973 35235 27031 35241
rect 28997 35275 29055 35281
rect 28997 35241 29009 35275
rect 29043 35272 29055 35275
rect 29270 35272 29276 35284
rect 29043 35244 29276 35272
rect 29043 35241 29055 35244
rect 28997 35235 29055 35241
rect 29270 35232 29276 35244
rect 29328 35232 29334 35284
rect 32493 35275 32551 35281
rect 32493 35241 32505 35275
rect 32539 35272 32551 35275
rect 32582 35272 32588 35284
rect 32539 35244 32588 35272
rect 32539 35241 32551 35244
rect 32493 35235 32551 35241
rect 32582 35232 32588 35244
rect 32640 35232 32646 35284
rect 42886 35272 42892 35284
rect 42847 35244 42892 35272
rect 42886 35232 42892 35244
rect 42944 35232 42950 35284
rect 44545 35275 44603 35281
rect 44545 35272 44557 35275
rect 43272 35244 44557 35272
rect 30101 35139 30159 35145
rect 30101 35136 30113 35139
rect 29196 35108 30113 35136
rect 24578 35028 24584 35080
rect 24636 35068 24642 35080
rect 29196 35077 29224 35108
rect 30101 35105 30113 35108
rect 30147 35105 30159 35139
rect 30558 35136 30564 35148
rect 30519 35108 30564 35136
rect 30101 35099 30159 35105
rect 30558 35096 30564 35108
rect 30616 35096 30622 35148
rect 33505 35139 33563 35145
rect 33505 35136 33517 35139
rect 32692 35108 33517 35136
rect 25593 35071 25651 35077
rect 25593 35068 25605 35071
rect 24636 35040 25605 35068
rect 24636 35028 24642 35040
rect 25593 35037 25605 35040
rect 25639 35037 25651 35071
rect 25593 35031 25651 35037
rect 25860 35071 25918 35077
rect 25860 35037 25872 35071
rect 25906 35037 25918 35071
rect 25860 35031 25918 35037
rect 29181 35071 29239 35077
rect 29181 35037 29193 35071
rect 29227 35037 29239 35071
rect 29181 35031 29239 35037
rect 29825 35071 29883 35077
rect 29825 35037 29837 35071
rect 29871 35037 29883 35071
rect 29825 35031 29883 35037
rect 29917 35071 29975 35077
rect 29917 35037 29929 35071
rect 29963 35068 29975 35071
rect 30466 35068 30472 35080
rect 29963 35040 30472 35068
rect 29963 35037 29975 35040
rect 29917 35031 29975 35037
rect 25608 34932 25636 35031
rect 25774 34960 25780 35012
rect 25832 35000 25838 35012
rect 25884 35000 25912 35031
rect 25832 34972 25912 35000
rect 29840 35000 29868 35031
rect 30466 35028 30472 35040
rect 30524 35068 30530 35080
rect 32692 35077 32720 35108
rect 33505 35105 33517 35108
rect 33551 35105 33563 35139
rect 40954 35136 40960 35148
rect 33505 35099 33563 35105
rect 40236 35108 40960 35136
rect 30745 35071 30803 35077
rect 30745 35068 30757 35071
rect 30524 35040 30757 35068
rect 30524 35028 30530 35040
rect 30745 35037 30757 35040
rect 30791 35037 30803 35071
rect 30745 35031 30803 35037
rect 30929 35071 30987 35077
rect 30929 35037 30941 35071
rect 30975 35068 30987 35071
rect 31573 35071 31631 35077
rect 31573 35068 31585 35071
rect 30975 35040 31585 35068
rect 30975 35037 30987 35040
rect 30929 35031 30987 35037
rect 31573 35037 31585 35040
rect 31619 35037 31631 35071
rect 31573 35031 31631 35037
rect 32677 35071 32735 35077
rect 32677 35037 32689 35071
rect 32723 35037 32735 35071
rect 33226 35068 33232 35080
rect 33187 35040 33232 35068
rect 32677 35031 32735 35037
rect 30374 35000 30380 35012
rect 29840 34972 30380 35000
rect 25832 34960 25838 34972
rect 30374 34960 30380 34972
rect 30432 34960 30438 35012
rect 30760 35000 30788 35031
rect 33226 35028 33232 35040
rect 33284 35028 33290 35080
rect 33321 35071 33379 35077
rect 33321 35037 33333 35071
rect 33367 35037 33379 35071
rect 33321 35031 33379 35037
rect 37829 35071 37887 35077
rect 37829 35037 37841 35071
rect 37875 35068 37887 35071
rect 38562 35068 38568 35080
rect 37875 35040 38568 35068
rect 37875 35037 37887 35040
rect 37829 35031 37887 35037
rect 33336 35000 33364 35031
rect 38562 35028 38568 35040
rect 38620 35028 38626 35080
rect 40236 35077 40264 35108
rect 40954 35096 40960 35108
rect 41012 35096 41018 35148
rect 40221 35071 40279 35077
rect 40221 35037 40233 35071
rect 40267 35037 40279 35071
rect 40402 35068 40408 35080
rect 40363 35040 40408 35068
rect 40221 35031 40279 35037
rect 40402 35028 40408 35040
rect 40460 35028 40466 35080
rect 40497 35071 40555 35077
rect 40497 35037 40509 35071
rect 40543 35068 40555 35071
rect 40678 35068 40684 35080
rect 40543 35040 40684 35068
rect 40543 35037 40555 35040
rect 40497 35031 40555 35037
rect 40678 35028 40684 35040
rect 40736 35028 40742 35080
rect 43162 35068 43168 35080
rect 43123 35040 43168 35068
rect 43162 35028 43168 35040
rect 43220 35028 43226 35080
rect 43272 35077 43300 35244
rect 44545 35241 44557 35244
rect 44591 35241 44603 35275
rect 44545 35235 44603 35241
rect 43346 35164 43352 35216
rect 43404 35204 43410 35216
rect 43404 35176 46980 35204
rect 43404 35164 43410 35176
rect 44269 35139 44327 35145
rect 44269 35105 44281 35139
rect 44315 35136 44327 35139
rect 44542 35136 44548 35148
rect 44315 35108 44548 35136
rect 44315 35105 44327 35108
rect 44269 35099 44327 35105
rect 44542 35096 44548 35108
rect 44600 35096 44606 35148
rect 45186 35096 45192 35148
rect 45244 35136 45250 35148
rect 45465 35139 45523 35145
rect 45465 35136 45477 35139
rect 45244 35108 45477 35136
rect 45244 35096 45250 35108
rect 45465 35105 45477 35108
rect 45511 35105 45523 35139
rect 45922 35136 45928 35148
rect 45883 35108 45928 35136
rect 45465 35099 45523 35105
rect 45922 35096 45928 35108
rect 45980 35096 45986 35148
rect 46952 35080 46980 35176
rect 43257 35071 43315 35077
rect 43257 35037 43269 35071
rect 43303 35037 43315 35071
rect 43257 35031 43315 35037
rect 43349 35071 43407 35077
rect 43349 35037 43361 35071
rect 43395 35068 43407 35071
rect 43438 35068 43444 35080
rect 43395 35040 43444 35068
rect 43395 35037 43407 35040
rect 43349 35031 43407 35037
rect 43438 35028 43444 35040
rect 43496 35028 43502 35080
rect 43530 35028 43536 35080
rect 43588 35068 43594 35080
rect 44174 35068 44180 35080
rect 43588 35040 43633 35068
rect 44135 35040 44180 35068
rect 43588 35028 43594 35040
rect 44174 35028 44180 35040
rect 44232 35028 44238 35080
rect 45557 35071 45615 35077
rect 45557 35037 45569 35071
rect 45603 35068 45615 35071
rect 46014 35068 46020 35080
rect 45603 35040 46020 35068
rect 45603 35037 45615 35040
rect 45557 35031 45615 35037
rect 46014 35028 46020 35040
rect 46072 35028 46078 35080
rect 46934 35068 46940 35080
rect 46895 35040 46940 35068
rect 46934 35028 46940 35040
rect 46992 35028 46998 35080
rect 47026 35028 47032 35080
rect 47084 35068 47090 35080
rect 47193 35071 47251 35077
rect 47193 35068 47205 35071
rect 47084 35040 47205 35068
rect 47084 35028 47090 35040
rect 47193 35037 47205 35040
rect 47239 35037 47251 35071
rect 47193 35031 47251 35037
rect 33870 35000 33876 35012
rect 30760 34972 33876 35000
rect 33870 34960 33876 34972
rect 33928 34960 33934 35012
rect 38841 35003 38899 35009
rect 38841 34969 38853 35003
rect 38887 35000 38899 35003
rect 39114 35000 39120 35012
rect 38887 34972 39120 35000
rect 38887 34969 38899 34972
rect 38841 34963 38899 34969
rect 39114 34960 39120 34972
rect 39172 34960 39178 35012
rect 42794 34960 42800 35012
rect 42852 35000 42858 35012
rect 43548 35000 43576 35028
rect 42852 34972 43576 35000
rect 42852 34960 42858 34972
rect 26050 34932 26056 34944
rect 25608 34904 26056 34932
rect 26050 34892 26056 34904
rect 26108 34892 26114 34944
rect 31386 34932 31392 34944
rect 31347 34904 31392 34932
rect 31386 34892 31392 34904
rect 31444 34892 31450 34944
rect 38010 34932 38016 34944
rect 37971 34904 38016 34932
rect 38010 34892 38016 34904
rect 38068 34892 38074 34944
rect 40037 34935 40095 34941
rect 40037 34901 40049 34935
rect 40083 34932 40095 34935
rect 40126 34932 40132 34944
rect 40083 34904 40132 34932
rect 40083 34901 40095 34904
rect 40037 34895 40095 34901
rect 40126 34892 40132 34904
rect 40184 34892 40190 34944
rect 46842 34892 46848 34944
rect 46900 34932 46906 34944
rect 48317 34935 48375 34941
rect 48317 34932 48329 34935
rect 46900 34904 48329 34932
rect 46900 34892 46906 34904
rect 48317 34901 48329 34904
rect 48363 34901 48375 34935
rect 48317 34895 48375 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 25314 34728 25320 34740
rect 25275 34700 25320 34728
rect 25314 34688 25320 34700
rect 25372 34688 25378 34740
rect 29641 34731 29699 34737
rect 29641 34697 29653 34731
rect 29687 34728 29699 34731
rect 30374 34728 30380 34740
rect 29687 34700 30380 34728
rect 29687 34697 29699 34700
rect 29641 34691 29699 34697
rect 30374 34688 30380 34700
rect 30432 34728 30438 34740
rect 31110 34728 31116 34740
rect 30432 34700 31116 34728
rect 30432 34688 30438 34700
rect 31110 34688 31116 34700
rect 31168 34688 31174 34740
rect 33226 34688 33232 34740
rect 33284 34728 33290 34740
rect 35434 34728 35440 34740
rect 33284 34700 35440 34728
rect 33284 34688 33290 34700
rect 35434 34688 35440 34700
rect 35492 34728 35498 34740
rect 35897 34731 35955 34737
rect 35897 34728 35909 34731
rect 35492 34700 35909 34728
rect 35492 34688 35498 34700
rect 35897 34697 35909 34700
rect 35943 34697 35955 34731
rect 39669 34731 39727 34737
rect 39669 34728 39681 34731
rect 35897 34691 35955 34697
rect 38764 34700 39681 34728
rect 24578 34660 24584 34672
rect 23952 34632 24584 34660
rect 23952 34601 23980 34632
rect 24578 34620 24584 34632
rect 24636 34620 24642 34672
rect 27522 34660 27528 34672
rect 27264 34632 27528 34660
rect 23937 34595 23995 34601
rect 23937 34561 23949 34595
rect 23983 34561 23995 34595
rect 23937 34555 23995 34561
rect 24026 34552 24032 34604
rect 24084 34592 24090 34604
rect 27264 34601 27292 34632
rect 27522 34620 27528 34632
rect 27580 34660 27586 34672
rect 29454 34660 29460 34672
rect 27580 34632 29460 34660
rect 27580 34620 27586 34632
rect 29454 34620 29460 34632
rect 29512 34620 29518 34672
rect 32122 34660 32128 34672
rect 30392 34632 32128 34660
rect 24193 34595 24251 34601
rect 24193 34592 24205 34595
rect 24084 34564 24205 34592
rect 24084 34552 24090 34564
rect 24193 34561 24205 34564
rect 24239 34561 24251 34595
rect 24193 34555 24251 34561
rect 27249 34595 27307 34601
rect 27249 34561 27261 34595
rect 27295 34561 27307 34595
rect 27249 34555 27307 34561
rect 27341 34595 27399 34601
rect 27341 34561 27353 34595
rect 27387 34592 27399 34595
rect 27430 34592 27436 34604
rect 27387 34564 27436 34592
rect 27387 34561 27399 34564
rect 27341 34555 27399 34561
rect 27430 34552 27436 34564
rect 27488 34552 27494 34604
rect 28074 34552 28080 34604
rect 28132 34592 28138 34604
rect 28261 34595 28319 34601
rect 28261 34592 28273 34595
rect 28132 34564 28273 34592
rect 28132 34552 28138 34564
rect 28261 34561 28273 34564
rect 28307 34561 28319 34595
rect 28261 34555 28319 34561
rect 28528 34595 28586 34601
rect 28528 34561 28540 34595
rect 28574 34592 28586 34595
rect 28902 34592 28908 34604
rect 28574 34564 28908 34592
rect 28574 34561 28586 34564
rect 28528 34555 28586 34561
rect 28902 34552 28908 34564
rect 28960 34552 28966 34604
rect 30392 34601 30420 34632
rect 32122 34620 32128 34632
rect 32180 34620 32186 34672
rect 38764 34604 38792 34700
rect 39669 34697 39681 34700
rect 39715 34697 39727 34731
rect 39669 34691 39727 34697
rect 43438 34688 43444 34740
rect 43496 34728 43502 34740
rect 43533 34731 43591 34737
rect 43533 34728 43545 34731
rect 43496 34700 43545 34728
rect 43496 34688 43502 34700
rect 43533 34697 43545 34700
rect 43579 34697 43591 34731
rect 43533 34691 43591 34697
rect 44174 34688 44180 34740
rect 44232 34728 44238 34740
rect 44453 34731 44511 34737
rect 44453 34728 44465 34731
rect 44232 34700 44465 34728
rect 44232 34688 44238 34700
rect 44453 34697 44465 34700
rect 44499 34697 44511 34731
rect 44453 34691 44511 34697
rect 46658 34688 46664 34740
rect 46716 34728 46722 34740
rect 47121 34731 47179 34737
rect 47121 34728 47133 34731
rect 46716 34700 47133 34728
rect 46716 34688 46722 34700
rect 47121 34697 47133 34700
rect 47167 34697 47179 34731
rect 47121 34691 47179 34697
rect 40034 34660 40040 34672
rect 39500 34632 40040 34660
rect 30377 34595 30435 34601
rect 30377 34561 30389 34595
rect 30423 34561 30435 34595
rect 30377 34555 30435 34561
rect 30644 34595 30702 34601
rect 30644 34561 30656 34595
rect 30690 34592 30702 34595
rect 31386 34592 31392 34604
rect 30690 34564 31392 34592
rect 30690 34561 30702 34564
rect 30644 34555 30702 34561
rect 31386 34552 31392 34564
rect 31444 34552 31450 34604
rect 33686 34592 33692 34604
rect 33647 34564 33692 34592
rect 33686 34552 33692 34564
rect 33744 34552 33750 34604
rect 33870 34592 33876 34604
rect 33831 34564 33876 34592
rect 33870 34552 33876 34564
rect 33928 34552 33934 34604
rect 34514 34592 34520 34604
rect 34475 34564 34520 34592
rect 34514 34552 34520 34564
rect 34572 34552 34578 34604
rect 34784 34595 34842 34601
rect 34784 34561 34796 34595
rect 34830 34592 34842 34595
rect 35710 34592 35716 34604
rect 34830 34564 35716 34592
rect 34830 34561 34842 34564
rect 34784 34555 34842 34561
rect 35710 34552 35716 34564
rect 35768 34552 35774 34604
rect 38197 34595 38255 34601
rect 38197 34561 38209 34595
rect 38243 34592 38255 34595
rect 38286 34592 38292 34604
rect 38243 34564 38292 34592
rect 38243 34561 38255 34564
rect 38197 34555 38255 34561
rect 38286 34552 38292 34564
rect 38344 34552 38350 34604
rect 38381 34595 38439 34601
rect 38381 34561 38393 34595
rect 38427 34592 38439 34595
rect 38746 34592 38752 34604
rect 38427 34564 38752 34592
rect 38427 34561 38439 34564
rect 38381 34555 38439 34561
rect 38746 34552 38752 34564
rect 38804 34552 38810 34604
rect 39500 34601 39528 34632
rect 40034 34620 40040 34632
rect 40092 34620 40098 34672
rect 40126 34620 40132 34672
rect 40184 34660 40190 34672
rect 40865 34663 40923 34669
rect 40865 34660 40877 34663
rect 40184 34632 40877 34660
rect 40184 34620 40190 34632
rect 40865 34629 40877 34632
rect 40911 34629 40923 34663
rect 40865 34623 40923 34629
rect 44085 34663 44143 34669
rect 44085 34629 44097 34663
rect 44131 34660 44143 34663
rect 44131 34632 45876 34660
rect 44131 34629 44143 34632
rect 44085 34623 44143 34629
rect 39485 34595 39543 34601
rect 39485 34561 39497 34595
rect 39531 34561 39543 34595
rect 39485 34555 39543 34561
rect 39761 34595 39819 34601
rect 39761 34561 39773 34595
rect 39807 34592 39819 34595
rect 40494 34592 40500 34604
rect 39807 34564 40500 34592
rect 39807 34561 39819 34564
rect 39761 34555 39819 34561
rect 40494 34552 40500 34564
rect 40552 34552 40558 34604
rect 43165 34595 43223 34601
rect 43165 34592 43177 34595
rect 41386 34564 43177 34592
rect 38565 34527 38623 34533
rect 38565 34493 38577 34527
rect 38611 34524 38623 34527
rect 38930 34524 38936 34536
rect 38611 34496 38936 34524
rect 38611 34493 38623 34496
rect 38565 34487 38623 34493
rect 38930 34484 38936 34496
rect 38988 34484 38994 34536
rect 39301 34527 39359 34533
rect 39301 34493 39313 34527
rect 39347 34524 39359 34527
rect 39390 34524 39396 34536
rect 39347 34496 39396 34524
rect 39347 34493 39359 34496
rect 39301 34487 39359 34493
rect 39390 34484 39396 34496
rect 39448 34484 39454 34536
rect 41386 34524 41414 34564
rect 43165 34561 43177 34564
rect 43211 34592 43223 34595
rect 43254 34592 43260 34604
rect 43211 34564 43260 34592
rect 43211 34561 43223 34564
rect 43165 34555 43223 34561
rect 43254 34552 43260 34564
rect 43312 34552 43318 34604
rect 43349 34595 43407 34601
rect 43349 34561 43361 34595
rect 43395 34561 43407 34595
rect 44266 34592 44272 34604
rect 44227 34564 44272 34592
rect 43349 34555 43407 34561
rect 39684 34496 41414 34524
rect 43364 34524 43392 34555
rect 44266 34552 44272 34564
rect 44324 34552 44330 34604
rect 44542 34592 44548 34604
rect 44503 34564 44548 34592
rect 44542 34552 44548 34564
rect 44600 34552 44606 34604
rect 45848 34601 45876 34632
rect 45833 34595 45891 34601
rect 45833 34561 45845 34595
rect 45879 34561 45891 34595
rect 45833 34555 45891 34561
rect 46014 34552 46020 34604
rect 46072 34592 46078 34604
rect 46842 34592 46848 34604
rect 46072 34564 46848 34592
rect 46072 34552 46078 34564
rect 46842 34552 46848 34564
rect 46900 34552 46906 34604
rect 44174 34524 44180 34536
rect 43364 34496 44180 34524
rect 38010 34416 38016 34468
rect 38068 34456 38074 34468
rect 38838 34456 38844 34468
rect 38068 34428 38844 34456
rect 38068 34416 38074 34428
rect 38838 34416 38844 34428
rect 38896 34456 38902 34468
rect 39684 34456 39712 34496
rect 44174 34484 44180 34496
rect 44232 34524 44238 34536
rect 44358 34524 44364 34536
rect 44232 34496 44364 34524
rect 44232 34484 44238 34496
rect 44358 34484 44364 34496
rect 44416 34484 44422 34536
rect 45922 34524 45928 34536
rect 45883 34496 45928 34524
rect 45922 34484 45928 34496
rect 45980 34484 45986 34536
rect 47121 34527 47179 34533
rect 47121 34493 47133 34527
rect 47167 34524 47179 34527
rect 47394 34524 47400 34536
rect 47167 34496 47400 34524
rect 47167 34493 47179 34496
rect 47121 34487 47179 34493
rect 47394 34484 47400 34496
rect 47452 34484 47458 34536
rect 41322 34456 41328 34468
rect 38896 34428 39712 34456
rect 40604 34428 41328 34456
rect 38896 34416 38902 34428
rect 27338 34348 27344 34400
rect 27396 34388 27402 34400
rect 27525 34391 27583 34397
rect 27525 34388 27537 34391
rect 27396 34360 27537 34388
rect 27396 34348 27402 34360
rect 27525 34357 27537 34360
rect 27571 34357 27583 34391
rect 27525 34351 27583 34357
rect 31754 34348 31760 34400
rect 31812 34388 31818 34400
rect 34057 34391 34115 34397
rect 31812 34360 31857 34388
rect 31812 34348 31818 34360
rect 34057 34357 34069 34391
rect 34103 34388 34115 34391
rect 34330 34388 34336 34400
rect 34103 34360 34336 34388
rect 34103 34357 34115 34360
rect 34057 34351 34115 34357
rect 34330 34348 34336 34360
rect 34388 34348 34394 34400
rect 37090 34348 37096 34400
rect 37148 34388 37154 34400
rect 40604 34388 40632 34428
rect 41322 34416 41328 34428
rect 41380 34416 41386 34468
rect 46201 34459 46259 34465
rect 46201 34425 46213 34459
rect 46247 34456 46259 34459
rect 47210 34456 47216 34468
rect 46247 34428 47216 34456
rect 46247 34425 46259 34428
rect 46201 34419 46259 34425
rect 47210 34416 47216 34428
rect 47268 34416 47274 34468
rect 37148 34360 40632 34388
rect 37148 34348 37154 34360
rect 40678 34348 40684 34400
rect 40736 34388 40742 34400
rect 40957 34391 41015 34397
rect 40957 34388 40969 34391
rect 40736 34360 40969 34388
rect 40736 34348 40742 34360
rect 40957 34357 40969 34360
rect 41003 34357 41015 34391
rect 40957 34351 41015 34357
rect 46937 34391 46995 34397
rect 46937 34357 46949 34391
rect 46983 34388 46995 34391
rect 47118 34388 47124 34400
rect 46983 34360 47124 34388
rect 46983 34357 46995 34360
rect 46937 34351 46995 34357
rect 47118 34348 47124 34360
rect 47176 34348 47182 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 28902 34184 28908 34196
rect 28863 34156 28908 34184
rect 28902 34144 28908 34156
rect 28960 34144 28966 34196
rect 35710 34184 35716 34196
rect 35671 34156 35716 34184
rect 35710 34144 35716 34156
rect 35768 34144 35774 34196
rect 43990 34184 43996 34196
rect 43951 34156 43996 34184
rect 43990 34144 43996 34156
rect 44048 34144 44054 34196
rect 48130 34184 48136 34196
rect 48091 34156 48136 34184
rect 48130 34144 48136 34156
rect 48188 34144 48194 34196
rect 33689 34119 33747 34125
rect 33689 34085 33701 34119
rect 33735 34116 33747 34119
rect 33870 34116 33876 34128
rect 33735 34088 33876 34116
rect 33735 34085 33747 34088
rect 33689 34079 33747 34085
rect 33870 34076 33876 34088
rect 33928 34076 33934 34128
rect 38105 34119 38163 34125
rect 38105 34085 38117 34119
rect 38151 34085 38163 34119
rect 38105 34079 38163 34085
rect 30101 34051 30159 34057
rect 30101 34048 30113 34051
rect 29104 34020 30113 34048
rect 26050 33980 26056 33992
rect 26011 33952 26056 33980
rect 26050 33940 26056 33952
rect 26108 33940 26114 33992
rect 29104 33989 29132 34020
rect 30101 34017 30113 34020
rect 30147 34017 30159 34051
rect 30101 34011 30159 34017
rect 34514 34008 34520 34060
rect 34572 34048 34578 34060
rect 36725 34051 36783 34057
rect 36725 34048 36737 34051
rect 34572 34020 36737 34048
rect 34572 34008 34578 34020
rect 36725 34017 36737 34020
rect 36771 34017 36783 34051
rect 36725 34011 36783 34017
rect 37734 34008 37740 34060
rect 37792 34048 37798 34060
rect 38120 34048 38148 34079
rect 38286 34076 38292 34128
rect 38344 34116 38350 34128
rect 40037 34119 40095 34125
rect 40037 34116 40049 34119
rect 38344 34088 40049 34116
rect 38344 34076 38350 34088
rect 40037 34085 40049 34088
rect 40083 34085 40095 34119
rect 40037 34079 40095 34085
rect 40773 34051 40831 34057
rect 40773 34048 40785 34051
rect 37792 34020 39620 34048
rect 37792 34008 37798 34020
rect 29089 33983 29147 33989
rect 29089 33949 29101 33983
rect 29135 33949 29147 33983
rect 29822 33980 29828 33992
rect 29783 33952 29828 33980
rect 29089 33943 29147 33949
rect 29822 33940 29828 33952
rect 29880 33940 29886 33992
rect 29917 33983 29975 33989
rect 29917 33949 29929 33983
rect 29963 33980 29975 33983
rect 30374 33980 30380 33992
rect 29963 33952 30380 33980
rect 29963 33949 29975 33952
rect 29917 33943 29975 33949
rect 30374 33940 30380 33952
rect 30432 33940 30438 33992
rect 30558 33940 30564 33992
rect 30616 33980 30622 33992
rect 31205 33983 31263 33989
rect 30616 33952 31064 33980
rect 30616 33940 30622 33952
rect 26320 33915 26378 33921
rect 26320 33881 26332 33915
rect 26366 33912 26378 33915
rect 27154 33912 27160 33924
rect 26366 33884 27160 33912
rect 26366 33881 26378 33884
rect 26320 33875 26378 33881
rect 27154 33872 27160 33884
rect 27212 33872 27218 33924
rect 29840 33912 29868 33940
rect 30929 33915 30987 33921
rect 30929 33912 30941 33915
rect 29840 33884 30941 33912
rect 30929 33881 30941 33884
rect 30975 33881 30987 33915
rect 31036 33912 31064 33952
rect 31205 33949 31217 33983
rect 31251 33980 31263 33983
rect 31754 33980 31760 33992
rect 31251 33952 31760 33980
rect 31251 33949 31263 33952
rect 31205 33943 31263 33949
rect 31754 33940 31760 33952
rect 31812 33940 31818 33992
rect 34330 33980 34336 33992
rect 34291 33952 34336 33980
rect 34330 33940 34336 33952
rect 34388 33940 34394 33992
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34848 33952 34897 33980
rect 34848 33940 34854 33952
rect 34885 33949 34897 33952
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 35069 33983 35127 33989
rect 35069 33949 35081 33983
rect 35115 33949 35127 33983
rect 35069 33943 35127 33949
rect 35253 33983 35311 33989
rect 35253 33949 35265 33983
rect 35299 33980 35311 33983
rect 35897 33983 35955 33989
rect 35897 33980 35909 33983
rect 35299 33952 35909 33980
rect 35299 33949 35311 33952
rect 35253 33943 35311 33949
rect 35897 33949 35909 33952
rect 35943 33949 35955 33983
rect 35897 33943 35955 33949
rect 38749 33983 38807 33989
rect 38749 33949 38761 33983
rect 38795 33949 38807 33983
rect 38930 33980 38936 33992
rect 38891 33952 38936 33980
rect 38749 33943 38807 33949
rect 31297 33915 31355 33921
rect 31297 33912 31309 33915
rect 31036 33884 31309 33912
rect 30929 33875 30987 33881
rect 31297 33881 31309 33884
rect 31343 33881 31355 33915
rect 33502 33912 33508 33924
rect 33463 33884 33508 33912
rect 31297 33875 31355 33881
rect 33502 33872 33508 33884
rect 33560 33872 33566 33924
rect 33870 33872 33876 33924
rect 33928 33912 33934 33924
rect 35084 33912 35112 33943
rect 33928 33884 35112 33912
rect 36992 33915 37050 33921
rect 33928 33872 33934 33884
rect 36992 33881 37004 33915
rect 37038 33912 37050 33915
rect 37458 33912 37464 33924
rect 37038 33884 37464 33912
rect 37038 33881 37050 33884
rect 36992 33875 37050 33881
rect 37458 33872 37464 33884
rect 37516 33872 37522 33924
rect 38764 33912 38792 33943
rect 38930 33940 38936 33952
rect 38988 33940 38994 33992
rect 39022 33940 39028 33992
rect 39080 33980 39086 33992
rect 39080 33952 39125 33980
rect 39080 33940 39086 33952
rect 39114 33912 39120 33924
rect 38764 33884 39120 33912
rect 39114 33872 39120 33884
rect 39172 33872 39178 33924
rect 39592 33912 39620 34020
rect 40236 34020 40785 34048
rect 40034 33980 40040 33992
rect 39995 33952 40040 33980
rect 40034 33940 40040 33952
rect 40092 33940 40098 33992
rect 40236 33989 40264 34020
rect 40773 34017 40785 34020
rect 40819 34017 40831 34051
rect 40773 34011 40831 34017
rect 40221 33983 40279 33989
rect 40221 33949 40233 33983
rect 40267 33949 40279 33983
rect 40678 33980 40684 33992
rect 40639 33952 40684 33980
rect 40221 33943 40279 33949
rect 40678 33940 40684 33952
rect 40736 33940 40742 33992
rect 40865 33983 40923 33989
rect 40865 33949 40877 33983
rect 40911 33980 40923 33983
rect 41046 33980 41052 33992
rect 40911 33952 41052 33980
rect 40911 33949 40923 33952
rect 40865 33943 40923 33949
rect 40494 33912 40500 33924
rect 39592 33884 40500 33912
rect 40494 33872 40500 33884
rect 40552 33912 40558 33924
rect 40880 33912 40908 33943
rect 41046 33940 41052 33952
rect 41104 33940 41110 33992
rect 43993 33983 44051 33989
rect 43993 33949 44005 33983
rect 44039 33949 44051 33983
rect 43993 33943 44051 33949
rect 40552 33884 40908 33912
rect 44008 33912 44036 33943
rect 44174 33940 44180 33992
rect 44232 33980 44238 33992
rect 45370 33980 45376 33992
rect 44232 33952 45376 33980
rect 44232 33940 44238 33952
rect 45370 33940 45376 33952
rect 45428 33940 45434 33992
rect 48314 33980 48320 33992
rect 48275 33952 48320 33980
rect 48314 33940 48320 33952
rect 48372 33940 48378 33992
rect 44008 33884 44220 33912
rect 40552 33872 40558 33884
rect 44192 33856 44220 33884
rect 27062 33804 27068 33856
rect 27120 33844 27126 33856
rect 27433 33847 27491 33853
rect 27433 33844 27445 33847
rect 27120 33816 27445 33844
rect 27120 33804 27126 33816
rect 27433 33813 27445 33816
rect 27479 33813 27491 33847
rect 31110 33844 31116 33856
rect 31071 33816 31116 33844
rect 27433 33807 27491 33813
rect 31110 33804 31116 33816
rect 31168 33804 31174 33856
rect 31481 33847 31539 33853
rect 31481 33813 31493 33847
rect 31527 33844 31539 33847
rect 32490 33844 32496 33856
rect 31527 33816 32496 33844
rect 31527 33813 31539 33816
rect 31481 33807 31539 33813
rect 32490 33804 32496 33816
rect 32548 33804 32554 33856
rect 34149 33847 34207 33853
rect 34149 33813 34161 33847
rect 34195 33844 34207 33847
rect 34514 33844 34520 33856
rect 34195 33816 34520 33844
rect 34195 33813 34207 33816
rect 34149 33807 34207 33813
rect 34514 33804 34520 33816
rect 34572 33804 34578 33856
rect 38194 33804 38200 33856
rect 38252 33844 38258 33856
rect 38565 33847 38623 33853
rect 38565 33844 38577 33847
rect 38252 33816 38577 33844
rect 38252 33804 38258 33816
rect 38565 33813 38577 33816
rect 38611 33813 38623 33847
rect 38565 33807 38623 33813
rect 44174 33804 44180 33856
rect 44232 33804 44238 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 27154 33640 27160 33652
rect 27115 33612 27160 33640
rect 27154 33600 27160 33612
rect 27212 33600 27218 33652
rect 27448 33612 34744 33640
rect 27448 33584 27476 33612
rect 25225 33575 25283 33581
rect 25225 33572 25237 33575
rect 24412 33544 25237 33572
rect 24412 33513 24440 33544
rect 25225 33541 25237 33544
rect 25271 33541 25283 33575
rect 27430 33572 27436 33584
rect 25225 33535 25283 33541
rect 27172 33544 27436 33572
rect 24397 33507 24455 33513
rect 24397 33473 24409 33507
rect 24443 33473 24455 33507
rect 24397 33467 24455 33473
rect 24946 33464 24952 33516
rect 25004 33504 25010 33516
rect 25041 33507 25099 33513
rect 25041 33504 25053 33507
rect 25004 33476 25053 33504
rect 25004 33464 25010 33476
rect 25041 33473 25053 33476
rect 25087 33504 25099 33507
rect 27172 33504 27200 33544
rect 27430 33532 27436 33544
rect 27488 33532 27494 33584
rect 30558 33532 30564 33584
rect 30616 33572 30622 33584
rect 30929 33575 30987 33581
rect 30929 33572 30941 33575
rect 30616 33544 30941 33572
rect 30616 33532 30622 33544
rect 30929 33541 30941 33544
rect 30975 33541 30987 33575
rect 30929 33535 30987 33541
rect 32122 33532 32128 33584
rect 32180 33572 32186 33584
rect 34514 33581 34520 33584
rect 34508 33572 34520 33581
rect 32180 33544 34284 33572
rect 34475 33544 34520 33572
rect 32180 33532 32186 33544
rect 27338 33504 27344 33516
rect 25087 33476 27200 33504
rect 27299 33476 27344 33504
rect 25087 33473 25099 33476
rect 25041 33467 25099 33473
rect 27338 33464 27344 33476
rect 27396 33464 27402 33516
rect 29822 33464 29828 33516
rect 29880 33504 29886 33516
rect 31205 33507 31263 33513
rect 31205 33504 31217 33507
rect 29880 33476 31217 33504
rect 29880 33464 29886 33476
rect 31205 33473 31217 33476
rect 31251 33473 31263 33507
rect 31205 33467 31263 33473
rect 33502 33464 33508 33516
rect 33560 33504 33566 33516
rect 34256 33513 34284 33544
rect 34508 33535 34520 33544
rect 34514 33532 34520 33535
rect 34572 33532 34578 33584
rect 34716 33572 34744 33612
rect 34790 33600 34796 33652
rect 34848 33640 34854 33652
rect 35621 33643 35679 33649
rect 35621 33640 35633 33643
rect 34848 33612 35633 33640
rect 34848 33600 34854 33612
rect 35621 33609 35633 33612
rect 35667 33609 35679 33643
rect 37458 33640 37464 33652
rect 37419 33612 37464 33640
rect 35621 33603 35679 33609
rect 37458 33600 37464 33612
rect 37516 33600 37522 33652
rect 38010 33640 38016 33652
rect 37844 33612 38016 33640
rect 36909 33575 36967 33581
rect 36909 33572 36921 33575
rect 34716 33544 36921 33572
rect 36909 33541 36921 33544
rect 36955 33572 36967 33575
rect 37090 33572 37096 33584
rect 36955 33544 37096 33572
rect 36955 33541 36967 33544
rect 36909 33535 36967 33541
rect 37090 33532 37096 33544
rect 37148 33532 37154 33584
rect 33597 33507 33655 33513
rect 33597 33504 33609 33507
rect 33560 33476 33609 33504
rect 33560 33464 33566 33476
rect 33597 33473 33609 33476
rect 33643 33473 33655 33507
rect 33597 33467 33655 33473
rect 34241 33507 34299 33513
rect 34241 33473 34253 33507
rect 34287 33473 34299 33507
rect 36541 33507 36599 33513
rect 36541 33504 36553 33507
rect 34241 33467 34299 33473
rect 34348 33476 36553 33504
rect 24857 33439 24915 33445
rect 24857 33405 24869 33439
rect 24903 33436 24915 33439
rect 26694 33436 26700 33448
rect 24903 33408 26700 33436
rect 24903 33405 24915 33408
rect 24857 33399 24915 33405
rect 26694 33396 26700 33408
rect 26752 33396 26758 33448
rect 31113 33439 31171 33445
rect 31113 33405 31125 33439
rect 31159 33436 31171 33439
rect 31754 33436 31760 33448
rect 31159 33408 31760 33436
rect 31159 33405 31171 33408
rect 31113 33399 31171 33405
rect 31754 33396 31760 33408
rect 31812 33396 31818 33448
rect 33410 33436 33416 33448
rect 33371 33408 33416 33436
rect 33410 33396 33416 33408
rect 33468 33396 33474 33448
rect 33612 33436 33640 33467
rect 34348 33436 34376 33476
rect 36541 33473 36553 33476
rect 36587 33504 36599 33507
rect 37550 33504 37556 33516
rect 36587 33476 37556 33504
rect 36587 33473 36599 33476
rect 36541 33467 36599 33473
rect 37550 33464 37556 33476
rect 37608 33464 37614 33516
rect 37734 33504 37740 33516
rect 37695 33476 37740 33504
rect 37734 33464 37740 33476
rect 37792 33464 37798 33516
rect 37844 33513 37872 33612
rect 38010 33600 38016 33612
rect 38068 33600 38074 33652
rect 38749 33643 38807 33649
rect 38749 33609 38761 33643
rect 38795 33640 38807 33643
rect 39022 33640 39028 33652
rect 38795 33612 39028 33640
rect 38795 33609 38807 33612
rect 38749 33603 38807 33609
rect 39022 33600 39028 33612
rect 39080 33600 39086 33652
rect 41414 33640 41420 33652
rect 39500 33612 41420 33640
rect 38194 33572 38200 33584
rect 37936 33544 38200 33572
rect 37936 33513 37964 33544
rect 38194 33532 38200 33544
rect 38252 33532 38258 33584
rect 37829 33507 37887 33513
rect 37829 33473 37841 33507
rect 37875 33473 37887 33507
rect 37829 33467 37887 33473
rect 37921 33507 37979 33513
rect 37921 33473 37933 33507
rect 37967 33473 37979 33507
rect 37921 33467 37979 33473
rect 38105 33507 38163 33513
rect 38105 33473 38117 33507
rect 38151 33473 38163 33507
rect 38105 33467 38163 33473
rect 33612 33408 34376 33436
rect 38120 33436 38148 33467
rect 38286 33464 38292 33516
rect 38344 33504 38350 33516
rect 38565 33507 38623 33513
rect 38565 33504 38577 33507
rect 38344 33476 38577 33504
rect 38344 33464 38350 33476
rect 38565 33473 38577 33476
rect 38611 33473 38623 33507
rect 38746 33504 38752 33516
rect 38707 33476 38752 33504
rect 38565 33467 38623 33473
rect 38746 33464 38752 33476
rect 38804 33464 38810 33516
rect 38930 33436 38936 33448
rect 38120 33408 38936 33436
rect 38930 33396 38936 33408
rect 38988 33436 38994 33448
rect 39500 33436 39528 33612
rect 41414 33600 41420 33612
rect 41472 33600 41478 33652
rect 40957 33575 41015 33581
rect 40957 33541 40969 33575
rect 41003 33572 41015 33575
rect 41230 33572 41236 33584
rect 41003 33544 41236 33572
rect 41003 33541 41015 33544
rect 40957 33535 41015 33541
rect 41230 33532 41236 33544
rect 41288 33532 41294 33584
rect 40773 33507 40831 33513
rect 40773 33473 40785 33507
rect 40819 33473 40831 33507
rect 40773 33467 40831 33473
rect 38988 33408 39528 33436
rect 40788 33436 40816 33467
rect 40862 33464 40868 33516
rect 40920 33504 40926 33516
rect 41049 33507 41107 33513
rect 41049 33504 41061 33507
rect 40920 33476 41061 33504
rect 40920 33464 40926 33476
rect 41049 33473 41061 33476
rect 41095 33473 41107 33507
rect 41049 33467 41107 33473
rect 45094 33464 45100 33516
rect 45152 33504 45158 33516
rect 45281 33507 45339 33513
rect 45281 33504 45293 33507
rect 45152 33476 45293 33504
rect 45152 33464 45158 33476
rect 45281 33473 45293 33476
rect 45327 33473 45339 33507
rect 45281 33467 45339 33473
rect 40788 33408 41092 33436
rect 38988 33396 38994 33408
rect 41064 33380 41092 33408
rect 44174 33396 44180 33448
rect 44232 33436 44238 33448
rect 45186 33436 45192 33448
rect 44232 33408 45192 33436
rect 44232 33396 44238 33408
rect 45186 33396 45192 33408
rect 45244 33396 45250 33448
rect 41046 33328 41052 33380
rect 41104 33328 41110 33380
rect 2314 33300 2320 33312
rect 2275 33272 2320 33300
rect 2314 33260 2320 33272
rect 2372 33260 2378 33312
rect 24213 33303 24271 33309
rect 24213 33269 24225 33303
rect 24259 33300 24271 33303
rect 24854 33300 24860 33312
rect 24259 33272 24860 33300
rect 24259 33269 24271 33272
rect 24213 33263 24271 33269
rect 24854 33260 24860 33272
rect 24912 33260 24918 33312
rect 31110 33300 31116 33312
rect 31071 33272 31116 33300
rect 31110 33260 31116 33272
rect 31168 33260 31174 33312
rect 31386 33300 31392 33312
rect 31347 33272 31392 33300
rect 31386 33260 31392 33272
rect 31444 33260 31450 33312
rect 33781 33303 33839 33309
rect 33781 33269 33793 33303
rect 33827 33300 33839 33303
rect 34146 33300 34152 33312
rect 33827 33272 34152 33300
rect 33827 33269 33839 33272
rect 33781 33263 33839 33269
rect 34146 33260 34152 33272
rect 34204 33260 34210 33312
rect 40773 33303 40831 33309
rect 40773 33269 40785 33303
rect 40819 33300 40831 33303
rect 41138 33300 41144 33312
rect 40819 33272 41144 33300
rect 40819 33269 40831 33272
rect 40773 33263 40831 33269
rect 41138 33260 41144 33272
rect 41196 33260 41202 33312
rect 45278 33260 45284 33312
rect 45336 33300 45342 33312
rect 45649 33303 45707 33309
rect 45649 33300 45661 33303
rect 45336 33272 45661 33300
rect 45336 33260 45342 33272
rect 45649 33269 45661 33272
rect 45695 33269 45707 33303
rect 47946 33300 47952 33312
rect 47907 33272 47952 33300
rect 45649 33263 45707 33269
rect 47946 33260 47952 33272
rect 48004 33260 48010 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 39114 33096 39120 33108
rect 39027 33068 39120 33096
rect 39114 33056 39120 33068
rect 39172 33096 39178 33108
rect 43162 33096 43168 33108
rect 39172 33068 43168 33096
rect 39172 33056 39178 33068
rect 43162 33056 43168 33068
rect 43220 33056 43226 33108
rect 44542 33056 44548 33108
rect 44600 33096 44606 33108
rect 45189 33099 45247 33105
rect 45189 33096 45201 33099
rect 44600 33068 45201 33096
rect 44600 33056 44606 33068
rect 45189 33065 45201 33068
rect 45235 33065 45247 33099
rect 45189 33059 45247 33065
rect 25958 32988 25964 33040
rect 26016 33028 26022 33040
rect 26694 33028 26700 33040
rect 26016 33000 26700 33028
rect 26016 32988 26022 33000
rect 26694 32988 26700 33000
rect 26752 32988 26758 33040
rect 1581 32963 1639 32969
rect 1581 32929 1593 32963
rect 1627 32960 1639 32963
rect 2314 32960 2320 32972
rect 1627 32932 2320 32960
rect 1627 32929 1639 32932
rect 1581 32923 1639 32929
rect 2314 32920 2320 32932
rect 2372 32920 2378 32972
rect 2774 32960 2780 32972
rect 2735 32932 2780 32960
rect 2774 32920 2780 32932
rect 2832 32920 2838 32972
rect 32122 32960 32128 32972
rect 32083 32932 32128 32960
rect 32122 32920 32128 32932
rect 32180 32920 32186 32972
rect 24581 32895 24639 32901
rect 24581 32861 24593 32895
rect 24627 32892 24639 32895
rect 26050 32892 26056 32904
rect 24627 32864 26056 32892
rect 24627 32861 24639 32864
rect 24581 32855 24639 32861
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 29917 32895 29975 32901
rect 29917 32861 29929 32895
rect 29963 32892 29975 32895
rect 30558 32892 30564 32904
rect 29963 32864 30564 32892
rect 29963 32861 29975 32864
rect 29917 32855 29975 32861
rect 30558 32852 30564 32864
rect 30616 32852 30622 32904
rect 31297 32895 31355 32901
rect 31297 32861 31309 32895
rect 31343 32892 31355 32895
rect 31386 32892 31392 32904
rect 31343 32864 31392 32892
rect 31343 32861 31355 32864
rect 31297 32855 31355 32861
rect 31386 32852 31392 32864
rect 31444 32852 31450 32904
rect 34146 32892 34152 32904
rect 34107 32864 34152 32892
rect 34146 32852 34152 32864
rect 34204 32852 34210 32904
rect 39132 32901 39160 33056
rect 44174 33028 44180 33040
rect 43456 33000 44180 33028
rect 40034 32920 40040 32972
rect 40092 32960 40098 32972
rect 40497 32963 40555 32969
rect 40497 32960 40509 32963
rect 40092 32932 40509 32960
rect 40092 32920 40098 32932
rect 40497 32929 40509 32932
rect 40543 32929 40555 32963
rect 40497 32923 40555 32929
rect 40957 32963 41015 32969
rect 40957 32929 40969 32963
rect 41003 32960 41015 32963
rect 41046 32960 41052 32972
rect 41003 32932 41052 32960
rect 41003 32929 41015 32932
rect 40957 32923 41015 32929
rect 41046 32920 41052 32932
rect 41104 32920 41110 32972
rect 42610 32920 42616 32972
rect 42668 32960 42674 32972
rect 43456 32969 43484 33000
rect 44174 32988 44180 33000
rect 44232 32988 44238 33040
rect 44284 33000 45508 33028
rect 43441 32963 43499 32969
rect 43441 32960 43453 32963
rect 42668 32932 43453 32960
rect 42668 32920 42674 32932
rect 43441 32929 43453 32932
rect 43487 32929 43499 32963
rect 43898 32960 43904 32972
rect 43811 32932 43904 32960
rect 43441 32923 43499 32929
rect 43898 32920 43904 32932
rect 43956 32960 43962 32972
rect 44284 32960 44312 33000
rect 43956 32932 44312 32960
rect 43956 32920 43962 32932
rect 36357 32895 36415 32901
rect 36357 32861 36369 32895
rect 36403 32892 36415 32895
rect 39117 32895 39175 32901
rect 36403 32864 37320 32892
rect 36403 32861 36415 32864
rect 36357 32855 36415 32861
rect 37292 32836 37320 32864
rect 39117 32861 39129 32895
rect 39163 32861 39175 32895
rect 39117 32855 39175 32861
rect 39393 32895 39451 32901
rect 39393 32861 39405 32895
rect 39439 32861 39451 32895
rect 39393 32855 39451 32861
rect 40589 32895 40647 32901
rect 40589 32861 40601 32895
rect 40635 32892 40647 32895
rect 41509 32895 41567 32901
rect 40635 32864 41414 32892
rect 40635 32861 40647 32864
rect 40589 32855 40647 32861
rect 1765 32827 1823 32833
rect 1765 32793 1777 32827
rect 1811 32824 1823 32827
rect 2406 32824 2412 32836
rect 1811 32796 2412 32824
rect 1811 32793 1823 32796
rect 1765 32787 1823 32793
rect 2406 32784 2412 32796
rect 2464 32784 2470 32836
rect 24854 32833 24860 32836
rect 24848 32824 24860 32833
rect 24815 32796 24860 32824
rect 24848 32787 24860 32796
rect 24854 32784 24860 32787
rect 24912 32784 24918 32836
rect 26418 32824 26424 32836
rect 26331 32796 26424 32824
rect 26418 32784 26424 32796
rect 26476 32824 26482 32836
rect 27522 32824 27528 32836
rect 26476 32796 27528 32824
rect 26476 32784 26482 32796
rect 27522 32784 27528 32796
rect 27580 32784 27586 32836
rect 31481 32827 31539 32833
rect 31481 32793 31493 32827
rect 31527 32824 31539 32827
rect 31754 32824 31760 32836
rect 31527 32796 31760 32824
rect 31527 32793 31539 32796
rect 31481 32787 31539 32793
rect 31754 32784 31760 32796
rect 31812 32784 31818 32836
rect 32398 32833 32404 32836
rect 32392 32787 32404 32833
rect 32456 32824 32462 32836
rect 36624 32827 36682 32833
rect 32456 32796 32492 32824
rect 32398 32784 32404 32787
rect 32456 32784 32462 32796
rect 36624 32793 36636 32827
rect 36670 32824 36682 32827
rect 37182 32824 37188 32836
rect 36670 32796 37188 32824
rect 36670 32793 36682 32796
rect 36624 32787 36682 32793
rect 37182 32784 37188 32796
rect 37240 32784 37246 32836
rect 37274 32784 37280 32836
rect 37332 32784 37338 32836
rect 39408 32824 39436 32855
rect 40862 32824 40868 32836
rect 39408 32796 40868 32824
rect 40862 32784 40868 32796
rect 40920 32784 40926 32836
rect 41386 32768 41414 32864
rect 41509 32861 41521 32895
rect 41555 32892 41567 32895
rect 43346 32892 43352 32904
rect 41555 32864 43352 32892
rect 41555 32861 41567 32864
rect 41509 32855 41567 32861
rect 43346 32852 43352 32864
rect 43404 32852 43410 32904
rect 43530 32892 43536 32904
rect 43491 32864 43536 32892
rect 43530 32852 43536 32864
rect 43588 32852 43594 32904
rect 44284 32902 44312 32932
rect 45278 32920 45284 32972
rect 45336 32960 45342 32972
rect 45480 32969 45508 33000
rect 45373 32963 45431 32969
rect 45373 32960 45385 32963
rect 45336 32932 45385 32960
rect 45336 32920 45342 32932
rect 45373 32929 45385 32932
rect 45419 32929 45431 32963
rect 45373 32923 45431 32929
rect 45465 32963 45523 32969
rect 45465 32929 45477 32963
rect 45511 32929 45523 32963
rect 45465 32923 45523 32929
rect 46477 32963 46535 32969
rect 46477 32929 46489 32963
rect 46523 32960 46535 32963
rect 47946 32960 47952 32972
rect 46523 32932 47952 32960
rect 46523 32929 46535 32932
rect 46477 32923 46535 32929
rect 47946 32920 47952 32932
rect 48004 32920 48010 32972
rect 44361 32905 44419 32911
rect 44361 32902 44373 32905
rect 44284 32874 44373 32902
rect 44361 32871 44373 32874
rect 44407 32871 44419 32905
rect 44542 32892 44548 32904
rect 44361 32865 44419 32871
rect 44503 32864 44548 32892
rect 44542 32852 44548 32864
rect 44600 32892 44606 32904
rect 45557 32895 45615 32901
rect 45388 32892 45509 32894
rect 45557 32892 45569 32895
rect 44600 32866 45569 32892
rect 44600 32864 45416 32866
rect 45481 32864 45569 32866
rect 44600 32852 44606 32864
rect 45557 32861 45569 32864
rect 45603 32861 45615 32895
rect 45557 32855 45615 32861
rect 45646 32852 45652 32904
rect 45704 32892 45710 32904
rect 45704 32864 45749 32892
rect 45704 32852 45710 32864
rect 41782 32833 41788 32836
rect 41776 32787 41788 32833
rect 41840 32824 41846 32836
rect 46661 32827 46719 32833
rect 41840 32796 41876 32824
rect 41782 32784 41788 32787
rect 41840 32784 41846 32796
rect 46661 32793 46673 32827
rect 46707 32824 46719 32827
rect 47854 32824 47860 32836
rect 46707 32796 47860 32824
rect 46707 32793 46719 32796
rect 46661 32787 46719 32793
rect 47854 32784 47860 32796
rect 47912 32784 47918 32836
rect 48314 32824 48320 32836
rect 48275 32796 48320 32824
rect 48314 32784 48320 32796
rect 48372 32784 48378 32836
rect 25961 32759 26019 32765
rect 25961 32725 25973 32759
rect 26007 32756 26019 32759
rect 26234 32756 26240 32768
rect 26007 32728 26240 32756
rect 26007 32725 26019 32728
rect 25961 32719 26019 32725
rect 26234 32716 26240 32728
rect 26292 32716 26298 32768
rect 26878 32756 26884 32768
rect 26839 32728 26884 32756
rect 26878 32716 26884 32728
rect 26936 32716 26942 32768
rect 29730 32756 29736 32768
rect 29691 32728 29736 32756
rect 29730 32716 29736 32728
rect 29788 32716 29794 32768
rect 31665 32759 31723 32765
rect 31665 32725 31677 32759
rect 31711 32756 31723 32759
rect 32766 32756 32772 32768
rect 31711 32728 32772 32756
rect 31711 32725 31723 32728
rect 31665 32719 31723 32725
rect 32766 32716 32772 32728
rect 32824 32716 32830 32768
rect 33410 32716 33416 32768
rect 33468 32756 33474 32768
rect 33505 32759 33563 32765
rect 33505 32756 33517 32759
rect 33468 32728 33517 32756
rect 33468 32716 33474 32728
rect 33505 32725 33517 32728
rect 33551 32725 33563 32759
rect 33962 32756 33968 32768
rect 33923 32728 33968 32756
rect 33505 32719 33563 32725
rect 33962 32716 33968 32728
rect 34020 32716 34026 32768
rect 37734 32756 37740 32768
rect 37695 32728 37740 32756
rect 37734 32716 37740 32728
rect 37792 32716 37798 32768
rect 38654 32716 38660 32768
rect 38712 32756 38718 32768
rect 38933 32759 38991 32765
rect 38933 32756 38945 32759
rect 38712 32728 38945 32756
rect 38712 32716 38718 32728
rect 38933 32725 38945 32728
rect 38979 32725 38991 32759
rect 38933 32719 38991 32725
rect 39301 32759 39359 32765
rect 39301 32725 39313 32759
rect 39347 32756 39359 32759
rect 40310 32756 40316 32768
rect 39347 32728 40316 32756
rect 39347 32725 39359 32728
rect 39301 32719 39359 32725
rect 40310 32716 40316 32728
rect 40368 32716 40374 32768
rect 41322 32716 41328 32768
rect 41380 32756 41414 32768
rect 42889 32759 42947 32765
rect 42889 32756 42901 32759
rect 41380 32728 42901 32756
rect 41380 32716 41386 32728
rect 42889 32725 42901 32728
rect 42935 32725 42947 32759
rect 42889 32719 42947 32725
rect 44545 32759 44603 32765
rect 44545 32725 44557 32759
rect 44591 32756 44603 32759
rect 44818 32756 44824 32768
rect 44591 32728 44824 32756
rect 44591 32725 44603 32728
rect 44545 32719 44603 32725
rect 44818 32716 44824 32728
rect 44876 32716 44882 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 2406 32552 2412 32564
rect 2367 32524 2412 32552
rect 2406 32512 2412 32524
rect 2464 32512 2470 32564
rect 26329 32555 26387 32561
rect 26329 32552 26341 32555
rect 25332 32524 26341 32552
rect 10502 32444 10508 32496
rect 10560 32484 10566 32496
rect 10560 32456 25268 32484
rect 10560 32444 10566 32456
rect 2317 32419 2375 32425
rect 2317 32385 2329 32419
rect 2363 32416 2375 32419
rect 2590 32416 2596 32428
rect 2363 32388 2596 32416
rect 2363 32385 2375 32388
rect 2317 32379 2375 32385
rect 2590 32376 2596 32388
rect 2648 32416 2654 32428
rect 7374 32416 7380 32428
rect 2648 32388 7380 32416
rect 2648 32376 2654 32388
rect 7374 32376 7380 32388
rect 7432 32376 7438 32428
rect 25133 32351 25191 32357
rect 25133 32317 25145 32351
rect 25179 32317 25191 32351
rect 25240 32348 25268 32456
rect 25332 32425 25360 32524
rect 26329 32521 26341 32524
rect 26375 32552 26387 32555
rect 27062 32552 27068 32564
rect 26375 32524 27068 32552
rect 26375 32521 26387 32524
rect 26329 32515 26387 32521
rect 27062 32512 27068 32524
rect 27120 32512 27126 32564
rect 29822 32512 29828 32564
rect 29880 32552 29886 32564
rect 30101 32555 30159 32561
rect 30101 32552 30113 32555
rect 29880 32524 30113 32552
rect 29880 32512 29886 32524
rect 30101 32521 30113 32524
rect 30147 32521 30159 32555
rect 30101 32515 30159 32521
rect 32309 32555 32367 32561
rect 32309 32521 32321 32555
rect 32355 32552 32367 32555
rect 32398 32552 32404 32564
rect 32355 32524 32404 32552
rect 32355 32521 32367 32524
rect 32309 32515 32367 32521
rect 32398 32512 32404 32524
rect 32456 32512 32462 32564
rect 32490 32512 32496 32564
rect 32548 32552 32554 32564
rect 41598 32552 41604 32564
rect 32548 32524 32628 32552
rect 32548 32512 32554 32524
rect 28988 32487 29046 32493
rect 25424 32456 28856 32484
rect 25317 32419 25375 32425
rect 25317 32385 25329 32419
rect 25363 32385 25375 32419
rect 25317 32379 25375 32385
rect 25424 32348 25452 32456
rect 25958 32416 25964 32428
rect 25919 32388 25964 32416
rect 25958 32376 25964 32388
rect 26016 32376 26022 32428
rect 26050 32376 26056 32428
rect 26108 32416 26114 32428
rect 28721 32419 28779 32425
rect 28721 32416 28733 32419
rect 26108 32388 28733 32416
rect 26108 32376 26114 32388
rect 28721 32385 28733 32388
rect 28767 32385 28779 32419
rect 28828 32416 28856 32456
rect 28988 32453 29000 32487
rect 29034 32484 29046 32487
rect 29730 32484 29736 32496
rect 29034 32456 29736 32484
rect 29034 32453 29046 32456
rect 28988 32447 29046 32453
rect 29730 32444 29736 32456
rect 29788 32444 29794 32496
rect 32600 32493 32628 32524
rect 36556 32524 41604 32552
rect 32585 32487 32643 32493
rect 32585 32453 32597 32487
rect 32631 32453 32643 32487
rect 32585 32447 32643 32453
rect 32766 32444 32772 32496
rect 32824 32493 32830 32496
rect 32824 32487 32853 32493
rect 32841 32453 32853 32487
rect 32824 32447 32853 32453
rect 32824 32444 32830 32447
rect 28828 32388 31754 32416
rect 28721 32379 28779 32385
rect 26234 32348 26240 32360
rect 25240 32320 25452 32348
rect 26147 32320 26240 32348
rect 25133 32311 25191 32317
rect 25148 32280 25176 32311
rect 26234 32308 26240 32320
rect 26292 32308 26298 32360
rect 26418 32308 26424 32360
rect 26476 32357 26482 32360
rect 26476 32351 26504 32357
rect 26492 32317 26504 32351
rect 26476 32311 26504 32317
rect 26476 32308 26482 32311
rect 26694 32308 26700 32360
rect 26752 32348 26758 32360
rect 27157 32351 27215 32357
rect 27157 32348 27169 32351
rect 26752 32320 27169 32348
rect 26752 32308 26758 32320
rect 27157 32317 27169 32320
rect 27203 32317 27215 32351
rect 27157 32311 27215 32317
rect 26252 32280 26280 32308
rect 27246 32280 27252 32292
rect 25148 32252 27252 32280
rect 27246 32240 27252 32252
rect 27304 32240 27310 32292
rect 27522 32280 27528 32292
rect 27483 32252 27528 32280
rect 27522 32240 27528 32252
rect 27580 32240 27586 32292
rect 31726 32280 31754 32388
rect 32398 32376 32404 32428
rect 32456 32416 32462 32428
rect 32493 32419 32551 32425
rect 32493 32416 32505 32419
rect 32456 32388 32505 32416
rect 32456 32376 32462 32388
rect 32493 32385 32505 32388
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 32677 32419 32735 32425
rect 32677 32385 32689 32419
rect 32723 32416 32735 32419
rect 32953 32419 33011 32425
rect 32723 32388 32812 32416
rect 32723 32385 32735 32388
rect 32677 32379 32735 32385
rect 32784 32360 32812 32388
rect 32953 32385 32965 32419
rect 32999 32416 33011 32419
rect 33962 32416 33968 32428
rect 32999 32388 33968 32416
rect 32999 32385 33011 32388
rect 32953 32379 33011 32385
rect 33962 32376 33968 32388
rect 34020 32376 34026 32428
rect 32766 32308 32772 32360
rect 32824 32348 32830 32360
rect 35526 32348 35532 32360
rect 32824 32320 35532 32348
rect 32824 32308 32830 32320
rect 35526 32308 35532 32320
rect 35584 32308 35590 32360
rect 36556 32280 36584 32524
rect 41598 32512 41604 32524
rect 41656 32512 41662 32564
rect 41693 32555 41751 32561
rect 41693 32521 41705 32555
rect 41739 32552 41751 32555
rect 41782 32552 41788 32564
rect 41739 32524 41788 32552
rect 41739 32521 41751 32524
rect 41693 32515 41751 32521
rect 41782 32512 41788 32524
rect 41840 32512 41846 32564
rect 41874 32512 41880 32564
rect 41932 32552 41938 32564
rect 43254 32552 43260 32564
rect 41932 32524 43260 32552
rect 41932 32512 41938 32524
rect 43254 32512 43260 32524
rect 43312 32512 43318 32564
rect 44818 32552 44824 32564
rect 44779 32524 44824 32552
rect 44818 32512 44824 32524
rect 44876 32512 44882 32564
rect 45278 32512 45284 32564
rect 45336 32552 45342 32564
rect 47854 32552 47860 32564
rect 45336 32524 46152 32552
rect 47815 32524 47860 32552
rect 45336 32512 45342 32524
rect 39114 32484 39120 32496
rect 37752 32456 39120 32484
rect 37458 32416 37464 32428
rect 37419 32388 37464 32416
rect 37458 32376 37464 32388
rect 37516 32376 37522 32428
rect 37550 32376 37556 32428
rect 37608 32416 37614 32428
rect 37752 32425 37780 32456
rect 39114 32444 39120 32456
rect 39172 32444 39178 32496
rect 41046 32484 41052 32496
rect 40696 32456 41052 32484
rect 37645 32419 37703 32425
rect 37645 32416 37657 32419
rect 37608 32388 37657 32416
rect 37608 32376 37614 32388
rect 37645 32385 37657 32388
rect 37691 32385 37703 32419
rect 37645 32379 37703 32385
rect 37737 32419 37795 32425
rect 37737 32385 37749 32419
rect 37783 32385 37795 32419
rect 37737 32379 37795 32385
rect 38933 32419 38991 32425
rect 38933 32385 38945 32419
rect 38979 32416 38991 32419
rect 39206 32416 39212 32428
rect 38979 32388 39212 32416
rect 38979 32385 38991 32388
rect 38933 32379 38991 32385
rect 39206 32376 39212 32388
rect 39264 32376 39270 32428
rect 40034 32416 40040 32428
rect 39500 32388 40040 32416
rect 39025 32351 39083 32357
rect 39025 32317 39037 32351
rect 39071 32348 39083 32351
rect 39500 32348 39528 32388
rect 40034 32376 40040 32388
rect 40092 32376 40098 32428
rect 40129 32419 40187 32425
rect 40129 32385 40141 32419
rect 40175 32414 40187 32419
rect 40696 32416 40724 32456
rect 41046 32444 41052 32456
rect 41104 32444 41110 32496
rect 41230 32444 41236 32496
rect 41288 32484 41294 32496
rect 42705 32487 42763 32493
rect 42705 32484 42717 32487
rect 41288 32456 42717 32484
rect 41288 32444 41294 32456
rect 42705 32453 42717 32456
rect 42751 32453 42763 32487
rect 42705 32447 42763 32453
rect 40957 32419 41015 32425
rect 40957 32416 40969 32419
rect 40236 32414 40724 32416
rect 40175 32388 40724 32414
rect 40788 32388 40969 32416
rect 40175 32386 40264 32388
rect 40175 32385 40187 32386
rect 40129 32379 40187 32385
rect 39071 32320 39528 32348
rect 40222 32351 40280 32357
rect 40222 32340 40234 32351
rect 39071 32317 39083 32320
rect 39025 32311 39083 32317
rect 40144 32317 40234 32340
rect 40268 32317 40280 32351
rect 40144 32312 40280 32317
rect 31726 32252 36584 32280
rect 37182 32240 37188 32292
rect 37240 32280 37246 32292
rect 37461 32283 37519 32289
rect 37461 32280 37473 32283
rect 37240 32252 37473 32280
rect 37240 32240 37246 32252
rect 37461 32249 37473 32252
rect 37507 32249 37519 32283
rect 37461 32243 37519 32249
rect 39301 32283 39359 32289
rect 39301 32249 39313 32283
rect 39347 32280 39359 32283
rect 40034 32280 40040 32292
rect 39347 32252 40040 32280
rect 39347 32249 39359 32252
rect 39301 32243 39359 32249
rect 40034 32240 40040 32252
rect 40092 32280 40098 32292
rect 40144 32280 40172 32312
rect 40222 32311 40280 32312
rect 40313 32351 40371 32357
rect 40313 32317 40325 32351
rect 40359 32317 40371 32351
rect 40313 32311 40371 32317
rect 40092 32252 40172 32280
rect 40328 32280 40356 32311
rect 40402 32308 40408 32360
rect 40460 32348 40466 32360
rect 40460 32320 40505 32348
rect 40460 32308 40466 32320
rect 40586 32280 40592 32292
rect 40328 32252 40592 32280
rect 40092 32240 40098 32252
rect 40586 32240 40592 32252
rect 40644 32240 40650 32292
rect 40788 32280 40816 32388
rect 40957 32385 40969 32388
rect 41003 32385 41015 32419
rect 41138 32416 41144 32428
rect 41099 32388 41144 32416
rect 40957 32379 41015 32385
rect 41138 32376 41144 32388
rect 41196 32376 41202 32428
rect 41414 32376 41420 32428
rect 41472 32416 41478 32428
rect 41509 32419 41567 32425
rect 41509 32416 41521 32419
rect 41472 32388 41521 32416
rect 41472 32376 41478 32388
rect 41509 32385 41521 32388
rect 41555 32385 41567 32419
rect 41509 32379 41567 32385
rect 41690 32376 41696 32428
rect 41748 32416 41754 32428
rect 42610 32416 42616 32428
rect 41748 32388 42616 32416
rect 41748 32376 41754 32388
rect 42610 32376 42616 32388
rect 42668 32376 42674 32428
rect 42797 32419 42855 32425
rect 42797 32385 42809 32419
rect 42843 32416 42855 32419
rect 42843 32388 42932 32416
rect 42843 32385 42855 32388
rect 42797 32379 42855 32385
rect 40862 32308 40868 32360
rect 40920 32348 40926 32360
rect 41233 32351 41291 32357
rect 41233 32348 41245 32351
rect 40920 32320 41245 32348
rect 40920 32308 40926 32320
rect 41233 32317 41245 32320
rect 41279 32317 41291 32351
rect 41233 32311 41291 32317
rect 41325 32351 41383 32357
rect 41325 32317 41337 32351
rect 41371 32348 41383 32351
rect 41874 32348 41880 32360
rect 41371 32320 41880 32348
rect 41371 32317 41383 32320
rect 41325 32311 41383 32317
rect 41874 32308 41880 32320
rect 41932 32308 41938 32360
rect 42702 32280 42708 32292
rect 40788 32252 42708 32280
rect 42702 32240 42708 32252
rect 42760 32240 42766 32292
rect 25501 32215 25559 32221
rect 25501 32181 25513 32215
rect 25547 32212 25559 32215
rect 26234 32212 26240 32224
rect 25547 32184 26240 32212
rect 25547 32181 25559 32184
rect 25501 32175 25559 32181
rect 26234 32172 26240 32184
rect 26292 32172 26298 32224
rect 26605 32215 26663 32221
rect 26605 32181 26617 32215
rect 26651 32212 26663 32215
rect 26786 32212 26792 32224
rect 26651 32184 26792 32212
rect 26651 32181 26663 32184
rect 26605 32175 26663 32181
rect 26786 32172 26792 32184
rect 26844 32172 26850 32224
rect 27614 32212 27620 32224
rect 27575 32184 27620 32212
rect 27614 32172 27620 32184
rect 27672 32172 27678 32224
rect 39945 32215 40003 32221
rect 39945 32181 39957 32215
rect 39991 32212 40003 32215
rect 40954 32212 40960 32224
rect 39991 32184 40960 32212
rect 39991 32181 40003 32184
rect 39945 32175 40003 32181
rect 40954 32172 40960 32184
rect 41012 32172 41018 32224
rect 41138 32172 41144 32224
rect 41196 32212 41202 32224
rect 42904 32212 42932 32388
rect 43162 32376 43168 32428
rect 43220 32416 43226 32428
rect 43625 32419 43683 32425
rect 43625 32416 43637 32419
rect 43220 32388 43637 32416
rect 43220 32376 43226 32388
rect 43625 32385 43637 32388
rect 43671 32385 43683 32419
rect 43806 32416 43812 32428
rect 43767 32388 43812 32416
rect 43625 32379 43683 32385
rect 43806 32376 43812 32388
rect 43864 32376 43870 32428
rect 43901 32419 43959 32425
rect 43901 32385 43913 32419
rect 43947 32416 43959 32419
rect 44836 32416 44864 32512
rect 45186 32444 45192 32496
rect 45244 32444 45250 32496
rect 43947 32388 44864 32416
rect 45204 32416 45232 32444
rect 46124 32425 46152 32524
rect 47854 32512 47860 32524
rect 47912 32512 47918 32564
rect 45281 32419 45339 32425
rect 45281 32416 45293 32419
rect 45204 32388 45293 32416
rect 43947 32385 43959 32388
rect 43901 32379 43959 32385
rect 45281 32385 45293 32388
rect 45327 32385 45339 32419
rect 45281 32379 45339 32385
rect 46109 32419 46167 32425
rect 46109 32385 46121 32419
rect 46155 32385 46167 32419
rect 46109 32379 46167 32385
rect 46658 32376 46664 32428
rect 46716 32416 46722 32428
rect 46937 32419 46995 32425
rect 46937 32416 46949 32419
rect 46716 32388 46949 32416
rect 46716 32376 46722 32388
rect 46937 32385 46949 32388
rect 46983 32385 46995 32419
rect 46937 32379 46995 32385
rect 47029 32419 47087 32425
rect 47029 32385 47041 32419
rect 47075 32416 47087 32419
rect 47118 32416 47124 32428
rect 47075 32388 47124 32416
rect 47075 32385 47087 32388
rect 47029 32379 47087 32385
rect 47118 32376 47124 32388
rect 47176 32376 47182 32428
rect 47765 32419 47823 32425
rect 47765 32385 47777 32419
rect 47811 32416 47823 32419
rect 47854 32416 47860 32428
rect 47811 32388 47860 32416
rect 47811 32385 47823 32388
rect 47765 32379 47823 32385
rect 47854 32376 47860 32388
rect 47912 32416 47918 32428
rect 48130 32416 48136 32428
rect 47912 32388 48136 32416
rect 47912 32376 47918 32388
rect 48130 32376 48136 32388
rect 48188 32376 48194 32428
rect 43530 32308 43536 32360
rect 43588 32348 43594 32360
rect 44082 32348 44088 32360
rect 43588 32320 44088 32348
rect 43588 32308 43594 32320
rect 44082 32308 44088 32320
rect 44140 32348 44146 32360
rect 45189 32351 45247 32357
rect 45189 32348 45201 32351
rect 44140 32320 45201 32348
rect 44140 32308 44146 32320
rect 45189 32317 45201 32320
rect 45235 32317 45247 32351
rect 45189 32311 45247 32317
rect 45465 32351 45523 32357
rect 45465 32317 45477 32351
rect 45511 32348 45523 32351
rect 46017 32351 46075 32357
rect 46017 32348 46029 32351
rect 45511 32320 46029 32348
rect 45511 32317 45523 32320
rect 45465 32311 45523 32317
rect 46017 32317 46029 32320
rect 46063 32317 46075 32351
rect 46017 32311 46075 32317
rect 47213 32351 47271 32357
rect 47213 32317 47225 32351
rect 47259 32348 47271 32351
rect 47394 32348 47400 32360
rect 47259 32320 47400 32348
rect 47259 32317 47271 32320
rect 47213 32311 47271 32317
rect 47394 32308 47400 32320
rect 47452 32308 47458 32360
rect 46474 32280 46480 32292
rect 46435 32252 46480 32280
rect 46474 32240 46480 32252
rect 46532 32240 46538 32292
rect 41196 32184 42932 32212
rect 41196 32172 41202 32184
rect 43346 32172 43352 32224
rect 43404 32212 43410 32224
rect 43441 32215 43499 32221
rect 43441 32212 43453 32215
rect 43404 32184 43453 32212
rect 43404 32172 43410 32184
rect 43441 32181 43453 32184
rect 43487 32181 43499 32215
rect 43441 32175 43499 32181
rect 47118 32172 47124 32224
rect 47176 32212 47182 32224
rect 47176 32184 47221 32212
rect 47176 32172 47182 32184
rect 47394 32172 47400 32224
rect 47452 32212 47458 32224
rect 47670 32212 47676 32224
rect 47452 32184 47676 32212
rect 47452 32172 47458 32184
rect 47670 32172 47676 32184
rect 47728 32172 47734 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 30558 32008 30564 32020
rect 30519 31980 30564 32008
rect 30558 31968 30564 31980
rect 30616 31968 30622 32020
rect 36722 31968 36728 32020
rect 36780 32008 36786 32020
rect 37182 32008 37188 32020
rect 36780 31980 37188 32008
rect 36780 31968 36786 31980
rect 37182 31968 37188 31980
rect 37240 32008 37246 32020
rect 37369 32011 37427 32017
rect 37369 32008 37381 32011
rect 37240 31980 37381 32008
rect 37240 31968 37246 31980
rect 37369 31977 37381 31980
rect 37415 31977 37427 32011
rect 37369 31971 37427 31977
rect 37458 31968 37464 32020
rect 37516 32008 37522 32020
rect 38289 32011 38347 32017
rect 38289 32008 38301 32011
rect 37516 31980 38301 32008
rect 37516 31968 37522 31980
rect 38289 31977 38301 31980
rect 38335 31977 38347 32011
rect 38289 31971 38347 31977
rect 39393 32011 39451 32017
rect 39393 31977 39405 32011
rect 39439 32008 39451 32011
rect 39439 31980 40264 32008
rect 39439 31977 39451 31980
rect 39393 31971 39451 31977
rect 26145 31943 26203 31949
rect 26145 31909 26157 31943
rect 26191 31940 26203 31943
rect 26326 31940 26332 31952
rect 26191 31912 26332 31940
rect 26191 31909 26203 31912
rect 26145 31903 26203 31909
rect 26326 31900 26332 31912
rect 26384 31900 26390 31952
rect 37090 31940 37096 31952
rect 34808 31912 37096 31940
rect 27157 31875 27215 31881
rect 27157 31872 27169 31875
rect 26620 31844 27169 31872
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31804 26387 31807
rect 26375 31776 26409 31804
rect 26375 31773 26387 31776
rect 26329 31767 26387 31773
rect 26344 31736 26372 31767
rect 26510 31764 26516 31816
rect 26568 31804 26574 31816
rect 26620 31813 26648 31844
rect 27157 31841 27169 31844
rect 27203 31841 27215 31875
rect 27157 31835 27215 31841
rect 26605 31807 26663 31813
rect 26605 31804 26617 31807
rect 26568 31776 26617 31804
rect 26568 31764 26574 31776
rect 26605 31773 26617 31776
rect 26651 31773 26663 31807
rect 27062 31804 27068 31816
rect 27023 31776 27068 31804
rect 26605 31767 26663 31773
rect 27062 31764 27068 31776
rect 27120 31764 27126 31816
rect 27246 31804 27252 31816
rect 27207 31776 27252 31804
rect 27246 31764 27252 31776
rect 27304 31764 27310 31816
rect 27801 31807 27859 31813
rect 27801 31773 27813 31807
rect 27847 31804 27859 31807
rect 29086 31804 29092 31816
rect 27847 31776 29092 31804
rect 27847 31773 27859 31776
rect 27801 31767 27859 31773
rect 29086 31764 29092 31776
rect 29144 31764 29150 31816
rect 30190 31804 30196 31816
rect 30151 31776 30196 31804
rect 30190 31764 30196 31776
rect 30248 31764 30254 31816
rect 30374 31804 30380 31816
rect 30335 31776 30380 31804
rect 30374 31764 30380 31776
rect 30432 31764 30438 31816
rect 34808 31804 34836 31912
rect 37090 31900 37096 31912
rect 37148 31900 37154 31952
rect 38746 31940 38752 31952
rect 38672 31912 38752 31940
rect 34885 31875 34943 31881
rect 34885 31841 34897 31875
rect 34931 31872 34943 31875
rect 35618 31872 35624 31884
rect 34931 31844 35624 31872
rect 34931 31841 34943 31844
rect 34885 31835 34943 31841
rect 35618 31832 35624 31844
rect 35676 31832 35682 31884
rect 37458 31832 37464 31884
rect 37516 31872 37522 31884
rect 37734 31872 37740 31884
rect 37516 31844 37740 31872
rect 37516 31832 37522 31844
rect 37734 31832 37740 31844
rect 37792 31872 37798 31884
rect 38672 31872 38700 31912
rect 38746 31900 38752 31912
rect 38804 31900 38810 31952
rect 40236 31940 40264 31980
rect 40310 31968 40316 32020
rect 40368 32008 40374 32020
rect 40405 32011 40463 32017
rect 40405 32008 40417 32011
rect 40368 31980 40417 32008
rect 40368 31968 40374 31980
rect 40405 31977 40417 31980
rect 40451 31977 40463 32011
rect 40862 32008 40868 32020
rect 40823 31980 40868 32008
rect 40405 31971 40463 31977
rect 40862 31968 40868 31980
rect 40920 31968 40926 32020
rect 43806 31968 43812 32020
rect 43864 32008 43870 32020
rect 44269 32011 44327 32017
rect 44269 32008 44281 32011
rect 43864 31980 44281 32008
rect 43864 31968 43870 31980
rect 44269 31977 44281 31980
rect 44315 31977 44327 32011
rect 44269 31971 44327 31977
rect 45189 32011 45247 32017
rect 45189 31977 45201 32011
rect 45235 32008 45247 32011
rect 45646 32008 45652 32020
rect 45235 31980 45652 32008
rect 45235 31977 45247 31980
rect 45189 31971 45247 31977
rect 45646 31968 45652 31980
rect 45704 31968 45710 32020
rect 46658 31968 46664 32020
rect 46716 32008 46722 32020
rect 48317 32011 48375 32017
rect 48317 32008 48329 32011
rect 46716 31980 48329 32008
rect 46716 31968 46722 31980
rect 48317 31977 48329 31980
rect 48363 31977 48375 32011
rect 48317 31971 48375 31977
rect 40770 31940 40776 31952
rect 40236 31912 40776 31940
rect 40770 31900 40776 31912
rect 40828 31900 40834 31952
rect 43162 31940 43168 31952
rect 41340 31912 43168 31940
rect 41046 31872 41052 31884
rect 37792 31844 38700 31872
rect 37792 31832 37798 31844
rect 35069 31807 35127 31813
rect 35069 31804 35081 31807
rect 34808 31776 35081 31804
rect 35069 31773 35081 31776
rect 35115 31773 35127 31807
rect 35069 31767 35127 31773
rect 35253 31807 35311 31813
rect 35253 31773 35265 31807
rect 35299 31804 35311 31807
rect 35894 31804 35900 31816
rect 35299 31776 35900 31804
rect 35299 31773 35311 31776
rect 35253 31767 35311 31773
rect 35894 31764 35900 31776
rect 35952 31764 35958 31816
rect 36078 31804 36084 31816
rect 36039 31776 36084 31804
rect 36078 31764 36084 31776
rect 36136 31764 36142 31816
rect 38378 31764 38384 31816
rect 38436 31804 38442 31816
rect 38672 31813 38700 31844
rect 39316 31844 40080 31872
rect 41007 31844 41052 31872
rect 38473 31807 38531 31813
rect 38473 31804 38485 31807
rect 38436 31776 38485 31804
rect 38436 31764 38442 31776
rect 38473 31773 38485 31776
rect 38519 31773 38531 31807
rect 38473 31767 38531 31773
rect 38657 31807 38715 31813
rect 38657 31773 38669 31807
rect 38703 31773 38715 31807
rect 38657 31767 38715 31773
rect 38749 31807 38807 31813
rect 38749 31773 38761 31807
rect 38795 31804 38807 31807
rect 38838 31804 38844 31816
rect 38795 31776 38844 31804
rect 38795 31773 38807 31776
rect 38749 31767 38807 31773
rect 26786 31736 26792 31748
rect 26344 31708 26792 31736
rect 26786 31696 26792 31708
rect 26844 31696 26850 31748
rect 26970 31696 26976 31748
rect 27028 31736 27034 31748
rect 28046 31739 28104 31745
rect 28046 31736 28058 31739
rect 27028 31708 28058 31736
rect 27028 31696 27034 31708
rect 28046 31705 28058 31708
rect 28092 31705 28104 31739
rect 28046 31699 28104 31705
rect 38562 31696 38568 31748
rect 38620 31736 38626 31748
rect 38764 31736 38792 31767
rect 38838 31764 38844 31776
rect 38896 31764 38902 31816
rect 39316 31813 39344 31844
rect 40052 31816 40080 31844
rect 41046 31832 41052 31844
rect 41104 31832 41110 31884
rect 41230 31872 41236 31884
rect 41191 31844 41236 31872
rect 41230 31832 41236 31844
rect 41288 31832 41294 31884
rect 41340 31881 41368 31912
rect 43162 31900 43168 31912
rect 43220 31900 43226 31952
rect 44082 31900 44088 31952
rect 44140 31940 44146 31952
rect 45557 31943 45615 31949
rect 45557 31940 45569 31943
rect 44140 31912 45569 31940
rect 44140 31900 44146 31912
rect 45557 31909 45569 31912
rect 45603 31909 45615 31943
rect 45557 31903 45615 31909
rect 41325 31875 41383 31881
rect 41325 31841 41337 31875
rect 41371 31841 41383 31875
rect 41325 31835 41383 31841
rect 45094 31832 45100 31884
rect 45152 31872 45158 31884
rect 45649 31875 45707 31881
rect 45649 31872 45661 31875
rect 45152 31844 45661 31872
rect 45152 31832 45158 31844
rect 45649 31841 45661 31844
rect 45695 31872 45707 31875
rect 46658 31872 46664 31884
rect 45695 31844 46664 31872
rect 45695 31841 45707 31844
rect 45649 31835 45707 31841
rect 46658 31832 46664 31844
rect 46716 31832 46722 31884
rect 46934 31872 46940 31884
rect 46895 31844 46940 31872
rect 46934 31832 46940 31844
rect 46992 31832 46998 31884
rect 39301 31807 39359 31813
rect 39301 31773 39313 31807
rect 39347 31773 39359 31807
rect 39301 31767 39359 31773
rect 39390 31764 39396 31816
rect 39448 31804 39454 31816
rect 39485 31807 39543 31813
rect 39485 31804 39497 31807
rect 39448 31776 39497 31804
rect 39448 31764 39454 31776
rect 39485 31773 39497 31776
rect 39531 31773 39543 31807
rect 40034 31804 40040 31816
rect 39995 31776 40040 31804
rect 39485 31767 39543 31773
rect 38620 31708 38792 31736
rect 39500 31736 39528 31767
rect 40034 31764 40040 31776
rect 40092 31764 40098 31816
rect 40586 31764 40592 31816
rect 40644 31764 40650 31816
rect 40770 31764 40776 31816
rect 40828 31804 40834 31816
rect 41141 31807 41199 31813
rect 41141 31804 41153 31807
rect 40828 31776 41153 31804
rect 40828 31764 40834 31776
rect 41141 31773 41153 31776
rect 41187 31773 41199 31807
rect 41141 31767 41199 31773
rect 43898 31764 43904 31816
rect 43956 31804 43962 31816
rect 43956 31776 44001 31804
rect 43956 31764 43962 31776
rect 45186 31764 45192 31816
rect 45244 31804 45250 31816
rect 45373 31807 45431 31813
rect 45373 31804 45385 31807
rect 45244 31776 45385 31804
rect 45244 31764 45250 31776
rect 45373 31773 45385 31776
rect 45419 31773 45431 31807
rect 45373 31767 45431 31773
rect 40221 31739 40279 31745
rect 40221 31736 40233 31739
rect 39500 31708 40233 31736
rect 38620 31696 38626 31708
rect 40221 31705 40233 31708
rect 40267 31736 40279 31739
rect 40604 31736 40632 31764
rect 40267 31708 40632 31736
rect 40267 31705 40279 31708
rect 40221 31699 40279 31705
rect 40954 31696 40960 31748
rect 41012 31736 41018 31748
rect 44085 31739 44143 31745
rect 44085 31736 44097 31739
rect 41012 31708 44097 31736
rect 41012 31696 41018 31708
rect 44085 31705 44097 31708
rect 44131 31736 44143 31739
rect 44542 31736 44548 31748
rect 44131 31708 44548 31736
rect 44131 31705 44143 31708
rect 44085 31699 44143 31705
rect 44542 31696 44548 31708
rect 44600 31696 44606 31748
rect 46934 31696 46940 31748
rect 46992 31736 46998 31748
rect 47182 31739 47240 31745
rect 47182 31736 47194 31739
rect 46992 31708 47194 31736
rect 46992 31696 46998 31708
rect 47182 31705 47194 31708
rect 47228 31705 47240 31739
rect 47182 31699 47240 31705
rect 26513 31671 26571 31677
rect 26513 31637 26525 31671
rect 26559 31668 26571 31671
rect 26602 31668 26608 31680
rect 26559 31640 26608 31668
rect 26559 31637 26571 31640
rect 26513 31631 26571 31637
rect 26602 31628 26608 31640
rect 26660 31668 26666 31680
rect 26878 31668 26884 31680
rect 26660 31640 26884 31668
rect 26660 31628 26666 31640
rect 26878 31628 26884 31640
rect 26936 31668 26942 31680
rect 27522 31668 27528 31680
rect 26936 31640 27528 31668
rect 26936 31628 26942 31640
rect 27522 31628 27528 31640
rect 27580 31628 27586 31680
rect 29181 31671 29239 31677
rect 29181 31637 29193 31671
rect 29227 31668 29239 31671
rect 29730 31668 29736 31680
rect 29227 31640 29736 31668
rect 29227 31637 29239 31640
rect 29181 31631 29239 31637
rect 29730 31628 29736 31640
rect 29788 31628 29794 31680
rect 39206 31628 39212 31680
rect 39264 31668 39270 31680
rect 40586 31668 40592 31680
rect 39264 31640 40592 31668
rect 39264 31628 39270 31640
rect 40586 31628 40592 31640
rect 40644 31628 40650 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 24857 31467 24915 31473
rect 24857 31433 24869 31467
rect 24903 31464 24915 31467
rect 26970 31464 26976 31476
rect 24903 31436 26976 31464
rect 24903 31433 24915 31436
rect 24857 31427 24915 31433
rect 26970 31424 26976 31436
rect 27028 31424 27034 31476
rect 28721 31467 28779 31473
rect 28721 31433 28733 31467
rect 28767 31433 28779 31467
rect 28721 31427 28779 31433
rect 24946 31396 24952 31408
rect 24136 31368 24952 31396
rect 24136 31337 24164 31368
rect 24946 31356 24952 31368
rect 25004 31356 25010 31408
rect 26528 31368 27384 31396
rect 26528 31340 26556 31368
rect 24121 31331 24179 31337
rect 24121 31297 24133 31331
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 24213 31331 24271 31337
rect 24213 31297 24225 31331
rect 24259 31328 24271 31331
rect 24302 31328 24308 31340
rect 24259 31300 24308 31328
rect 24259 31297 24271 31300
rect 24213 31291 24271 31297
rect 24302 31288 24308 31300
rect 24360 31288 24366 31340
rect 24397 31331 24455 31337
rect 24397 31297 24409 31331
rect 24443 31328 24455 31331
rect 25041 31331 25099 31337
rect 25041 31328 25053 31331
rect 24443 31300 25053 31328
rect 24443 31297 24455 31300
rect 24397 31291 24455 31297
rect 25041 31297 25053 31300
rect 25087 31297 25099 31331
rect 26234 31328 26240 31340
rect 26147 31300 26240 31328
rect 25041 31291 25099 31297
rect 26234 31288 26240 31300
rect 26292 31288 26298 31340
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31328 26387 31331
rect 26510 31328 26516 31340
rect 26375 31300 26516 31328
rect 26375 31297 26387 31300
rect 26329 31291 26387 31297
rect 26510 31288 26516 31300
rect 26568 31288 26574 31340
rect 27154 31328 27160 31340
rect 27115 31300 27160 31328
rect 27154 31288 27160 31300
rect 27212 31288 27218 31340
rect 27356 31337 27384 31368
rect 27522 31356 27528 31408
rect 27580 31396 27586 31408
rect 28736 31396 28764 31427
rect 29730 31424 29736 31476
rect 29788 31464 29794 31476
rect 29788 31436 31616 31464
rect 29788 31424 29794 31436
rect 29610 31399 29668 31405
rect 29610 31396 29622 31399
rect 27580 31368 27752 31396
rect 28736 31368 29622 31396
rect 27580 31356 27586 31368
rect 27341 31331 27399 31337
rect 27341 31297 27353 31331
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 27433 31331 27491 31337
rect 27433 31297 27445 31331
rect 27479 31328 27491 31331
rect 27614 31328 27620 31340
rect 27479 31300 27620 31328
rect 27479 31297 27491 31300
rect 27433 31291 27491 31297
rect 26050 31124 26056 31136
rect 26011 31096 26056 31124
rect 26050 31084 26056 31096
rect 26108 31084 26114 31136
rect 26252 31124 26280 31288
rect 26602 31260 26608 31272
rect 26563 31232 26608 31260
rect 26602 31220 26608 31232
rect 26660 31220 26666 31272
rect 26513 31195 26571 31201
rect 26513 31161 26525 31195
rect 26559 31192 26571 31195
rect 27448 31192 27476 31291
rect 27614 31288 27620 31300
rect 27672 31288 27678 31340
rect 27724 31337 27752 31368
rect 29610 31365 29622 31368
rect 29656 31365 29668 31399
rect 29610 31359 29668 31365
rect 30190 31356 30196 31408
rect 30248 31396 30254 31408
rect 31297 31399 31355 31405
rect 31297 31396 31309 31399
rect 30248 31368 31309 31396
rect 30248 31356 30254 31368
rect 31297 31365 31309 31368
rect 31343 31365 31355 31399
rect 31297 31359 31355 31365
rect 27709 31331 27767 31337
rect 27709 31297 27721 31331
rect 27755 31297 27767 31331
rect 27709 31291 27767 31297
rect 28905 31331 28963 31337
rect 28905 31297 28917 31331
rect 28951 31328 28963 31331
rect 30098 31328 30104 31340
rect 28951 31300 30104 31328
rect 28951 31297 28963 31300
rect 28905 31291 28963 31297
rect 30098 31288 30104 31300
rect 30156 31288 30162 31340
rect 27525 31263 27583 31269
rect 27525 31229 27537 31263
rect 27571 31229 27583 31263
rect 27525 31223 27583 31229
rect 26559 31164 27476 31192
rect 26559 31161 26571 31164
rect 26513 31155 26571 31161
rect 27540 31124 27568 31223
rect 29086 31220 29092 31272
rect 29144 31260 29150 31272
rect 29362 31260 29368 31272
rect 29144 31232 29368 31260
rect 29144 31220 29150 31232
rect 29362 31220 29368 31232
rect 29420 31220 29426 31272
rect 31312 31192 31340 31359
rect 31588 31337 31616 31436
rect 31754 31424 31760 31476
rect 31812 31464 31818 31476
rect 31812 31436 31857 31464
rect 31812 31424 31818 31436
rect 32398 31424 32404 31476
rect 32456 31464 32462 31476
rect 32861 31467 32919 31473
rect 32861 31464 32873 31467
rect 32456 31436 32873 31464
rect 32456 31424 32462 31436
rect 32861 31433 32873 31436
rect 32907 31433 32919 31467
rect 37550 31464 37556 31476
rect 37511 31436 37556 31464
rect 32861 31427 32919 31433
rect 37550 31424 37556 31436
rect 37608 31464 37614 31476
rect 38838 31464 38844 31476
rect 37608 31436 38844 31464
rect 37608 31424 37614 31436
rect 38838 31424 38844 31436
rect 38896 31424 38902 31476
rect 40402 31424 40408 31476
rect 40460 31464 40466 31476
rect 40773 31467 40831 31473
rect 40773 31464 40785 31467
rect 40460 31436 40785 31464
rect 40460 31424 40466 31436
rect 40773 31433 40785 31436
rect 40819 31433 40831 31467
rect 47026 31464 47032 31476
rect 46987 31436 47032 31464
rect 40773 31427 40831 31433
rect 47026 31424 47032 31436
rect 47084 31424 47090 31476
rect 47118 31424 47124 31476
rect 47176 31424 47182 31476
rect 32122 31356 32128 31408
rect 32180 31396 32186 31408
rect 32585 31399 32643 31405
rect 32585 31396 32597 31399
rect 32180 31368 32597 31396
rect 32180 31356 32186 31368
rect 32585 31365 32597 31368
rect 32631 31365 32643 31399
rect 32585 31359 32643 31365
rect 33962 31356 33968 31408
rect 34020 31396 34026 31408
rect 34302 31399 34360 31405
rect 34302 31396 34314 31399
rect 34020 31368 34314 31396
rect 34020 31356 34026 31368
rect 34302 31365 34314 31368
rect 34348 31365 34360 31399
rect 39206 31396 39212 31408
rect 34302 31359 34360 31365
rect 38396 31368 39212 31396
rect 31573 31331 31631 31337
rect 31573 31297 31585 31331
rect 31619 31328 31631 31331
rect 32309 31331 32367 31337
rect 32309 31328 32321 31331
rect 31619 31300 32321 31328
rect 31619 31297 31631 31300
rect 31573 31291 31631 31297
rect 32309 31297 32321 31300
rect 32355 31297 32367 31331
rect 32490 31328 32496 31340
rect 32451 31300 32496 31328
rect 32309 31291 32367 31297
rect 32490 31288 32496 31300
rect 32548 31288 32554 31340
rect 32677 31331 32735 31337
rect 32677 31297 32689 31331
rect 32723 31297 32735 31331
rect 32677 31291 32735 31297
rect 31481 31263 31539 31269
rect 31481 31229 31493 31263
rect 31527 31260 31539 31263
rect 32122 31260 32128 31272
rect 31527 31232 32128 31260
rect 31527 31229 31539 31232
rect 31481 31223 31539 31229
rect 32122 31220 32128 31232
rect 32180 31220 32186 31272
rect 32692 31192 32720 31291
rect 35894 31288 35900 31340
rect 35952 31328 35958 31340
rect 36081 31331 36139 31337
rect 36081 31328 36093 31331
rect 35952 31300 36093 31328
rect 35952 31288 35958 31300
rect 36081 31297 36093 31300
rect 36127 31297 36139 31331
rect 37458 31328 37464 31340
rect 37419 31300 37464 31328
rect 36081 31291 36139 31297
rect 37458 31288 37464 31300
rect 37516 31288 37522 31340
rect 38396 31337 38424 31368
rect 39206 31356 39212 31368
rect 39264 31356 39270 31408
rect 46845 31399 46903 31405
rect 46845 31365 46857 31399
rect 46891 31396 46903 31399
rect 47136 31396 47164 31424
rect 46891 31368 47164 31396
rect 46891 31365 46903 31368
rect 46845 31359 46903 31365
rect 38381 31331 38439 31337
rect 38381 31297 38393 31331
rect 38427 31297 38439 31331
rect 38381 31291 38439 31297
rect 38473 31331 38531 31337
rect 38473 31297 38485 31331
rect 38519 31297 38531 31331
rect 38473 31291 38531 31297
rect 38565 31331 38623 31337
rect 38565 31297 38577 31331
rect 38611 31328 38623 31331
rect 38654 31328 38660 31340
rect 38611 31300 38660 31328
rect 38611 31297 38623 31300
rect 38565 31291 38623 31297
rect 34054 31260 34060 31272
rect 34015 31232 34060 31260
rect 34054 31220 34060 31232
rect 34112 31220 34118 31272
rect 33594 31192 33600 31204
rect 31312 31164 33600 31192
rect 33594 31152 33600 31164
rect 33652 31152 33658 31204
rect 38488 31192 38516 31291
rect 38654 31288 38660 31300
rect 38712 31288 38718 31340
rect 38746 31288 38752 31340
rect 38804 31328 38810 31340
rect 38930 31328 38936 31340
rect 38804 31300 38936 31328
rect 38804 31288 38810 31300
rect 38930 31288 38936 31300
rect 38988 31288 38994 31340
rect 40678 31288 40684 31340
rect 40736 31328 40742 31340
rect 40957 31331 41015 31337
rect 40957 31328 40969 31331
rect 40736 31300 40969 31328
rect 40736 31288 40742 31300
rect 40957 31297 40969 31300
rect 41003 31328 41015 31331
rect 41598 31328 41604 31340
rect 41003 31300 41604 31328
rect 41003 31297 41015 31300
rect 40957 31291 41015 31297
rect 41598 31288 41604 31300
rect 41656 31288 41662 31340
rect 46474 31288 46480 31340
rect 46532 31328 46538 31340
rect 47121 31331 47179 31337
rect 47121 31328 47133 31331
rect 46532 31300 47133 31328
rect 46532 31288 46538 31300
rect 47121 31297 47133 31300
rect 47167 31297 47179 31331
rect 47121 31291 47179 31297
rect 40586 31220 40592 31272
rect 40644 31260 40650 31272
rect 41138 31260 41144 31272
rect 40644 31232 41144 31260
rect 40644 31220 40650 31232
rect 41138 31220 41144 31232
rect 41196 31220 41202 31272
rect 41233 31263 41291 31269
rect 41233 31229 41245 31263
rect 41279 31260 41291 31263
rect 41322 31260 41328 31272
rect 41279 31232 41328 31260
rect 41279 31229 41291 31232
rect 41233 31223 41291 31229
rect 41322 31220 41328 31232
rect 41380 31220 41386 31272
rect 42794 31220 42800 31272
rect 42852 31260 42858 31272
rect 43530 31260 43536 31272
rect 42852 31232 43536 31260
rect 42852 31220 42858 31232
rect 43530 31220 43536 31232
rect 43588 31220 43594 31272
rect 38562 31192 38568 31204
rect 38488 31164 38568 31192
rect 38562 31152 38568 31164
rect 38620 31152 38626 31204
rect 46845 31195 46903 31201
rect 46845 31161 46857 31195
rect 46891 31192 46903 31195
rect 46934 31192 46940 31204
rect 46891 31164 46940 31192
rect 46891 31161 46903 31164
rect 46845 31155 46903 31161
rect 46934 31152 46940 31164
rect 46992 31152 46998 31204
rect 27890 31124 27896 31136
rect 26252 31096 27568 31124
rect 27851 31096 27896 31124
rect 27890 31084 27896 31096
rect 27948 31084 27954 31136
rect 30745 31127 30803 31133
rect 30745 31093 30757 31127
rect 30791 31124 30803 31127
rect 31202 31124 31208 31136
rect 30791 31096 31208 31124
rect 30791 31093 30803 31096
rect 30745 31087 30803 31093
rect 31202 31084 31208 31096
rect 31260 31124 31266 31136
rect 31573 31127 31631 31133
rect 31573 31124 31585 31127
rect 31260 31096 31585 31124
rect 31260 31084 31266 31096
rect 31573 31093 31585 31096
rect 31619 31124 31631 31127
rect 32490 31124 32496 31136
rect 31619 31096 32496 31124
rect 31619 31093 31631 31096
rect 31573 31087 31631 31093
rect 32490 31084 32496 31096
rect 32548 31084 32554 31136
rect 35434 31124 35440 31136
rect 35395 31096 35440 31124
rect 35434 31084 35440 31096
rect 35492 31084 35498 31136
rect 35894 31124 35900 31136
rect 35855 31096 35900 31124
rect 35894 31084 35900 31096
rect 35952 31084 35958 31136
rect 38102 31124 38108 31136
rect 38063 31096 38108 31124
rect 38102 31084 38108 31096
rect 38160 31084 38166 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 30098 30920 30104 30932
rect 30059 30892 30104 30920
rect 30098 30880 30104 30892
rect 30156 30880 30162 30932
rect 33594 30920 33600 30932
rect 33555 30892 33600 30920
rect 33594 30880 33600 30892
rect 33652 30880 33658 30932
rect 38841 30923 38899 30929
rect 38841 30889 38853 30923
rect 38887 30920 38899 30923
rect 40586 30920 40592 30932
rect 38887 30892 40592 30920
rect 38887 30889 38899 30892
rect 38841 30883 38899 30889
rect 40586 30880 40592 30892
rect 40644 30880 40650 30932
rect 44082 30920 44088 30932
rect 43272 30892 44088 30920
rect 29730 30784 29736 30796
rect 29691 30756 29736 30784
rect 29730 30744 29736 30756
rect 29788 30744 29794 30796
rect 31202 30784 31208 30796
rect 31163 30756 31208 30784
rect 31202 30744 31208 30756
rect 31260 30744 31266 30796
rect 40313 30787 40371 30793
rect 40313 30753 40325 30787
rect 40359 30784 40371 30787
rect 42334 30784 42340 30796
rect 40359 30756 42340 30784
rect 40359 30753 40371 30756
rect 40313 30747 40371 30753
rect 42334 30744 42340 30756
rect 42392 30744 42398 30796
rect 43272 30784 43300 30892
rect 44082 30880 44088 30892
rect 44140 30880 44146 30932
rect 45830 30920 45836 30932
rect 45791 30892 45836 30920
rect 45830 30880 45836 30892
rect 45888 30880 45894 30932
rect 43346 30812 43352 30864
rect 43404 30812 43410 30864
rect 43180 30756 43300 30784
rect 26510 30716 26516 30728
rect 26471 30688 26516 30716
rect 26510 30676 26516 30688
rect 26568 30676 26574 30728
rect 26602 30676 26608 30728
rect 26660 30716 26666 30728
rect 26786 30716 26792 30728
rect 26660 30688 26705 30716
rect 26747 30688 26792 30716
rect 26660 30676 26666 30688
rect 26786 30676 26792 30688
rect 26844 30676 26850 30728
rect 26881 30719 26939 30725
rect 26881 30685 26893 30719
rect 26927 30716 26939 30719
rect 27154 30716 27160 30728
rect 26927 30688 27160 30716
rect 26927 30685 26939 30688
rect 26881 30679 26939 30685
rect 27154 30676 27160 30688
rect 27212 30716 27218 30728
rect 27430 30716 27436 30728
rect 27212 30688 27436 30716
rect 27212 30676 27218 30688
rect 27430 30676 27436 30688
rect 27488 30676 27494 30728
rect 29917 30719 29975 30725
rect 29917 30685 29929 30719
rect 29963 30716 29975 30719
rect 30374 30716 30380 30728
rect 29963 30688 30380 30716
rect 29963 30685 29975 30688
rect 29917 30679 29975 30685
rect 30374 30676 30380 30688
rect 30432 30716 30438 30728
rect 31386 30716 31392 30728
rect 30432 30688 31392 30716
rect 30432 30676 30438 30688
rect 31386 30676 31392 30688
rect 31444 30676 31450 30728
rect 32214 30716 32220 30728
rect 32175 30688 32220 30716
rect 32214 30676 32220 30688
rect 32272 30676 32278 30728
rect 34054 30676 34060 30728
rect 34112 30716 34118 30728
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 34112 30688 34897 30716
rect 34112 30676 34118 30688
rect 34885 30685 34897 30688
rect 34931 30716 34943 30719
rect 37458 30716 37464 30728
rect 34931 30688 37464 30716
rect 34931 30685 34943 30688
rect 34885 30679 34943 30685
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 37728 30719 37786 30725
rect 37728 30685 37740 30719
rect 37774 30716 37786 30719
rect 38102 30716 38108 30728
rect 37774 30688 38108 30716
rect 37774 30685 37786 30688
rect 37728 30679 37786 30685
rect 38102 30676 38108 30688
rect 38160 30676 38166 30728
rect 40497 30719 40555 30725
rect 40497 30685 40509 30719
rect 40543 30685 40555 30719
rect 40770 30716 40776 30728
rect 40731 30688 40776 30716
rect 40497 30679 40555 30685
rect 32484 30651 32542 30657
rect 32484 30617 32496 30651
rect 32530 30648 32542 30651
rect 33134 30648 33140 30660
rect 32530 30620 33140 30648
rect 32530 30617 32542 30620
rect 32484 30611 32542 30617
rect 33134 30608 33140 30620
rect 33192 30608 33198 30660
rect 35152 30651 35210 30657
rect 35152 30617 35164 30651
rect 35198 30648 35210 30651
rect 35894 30648 35900 30660
rect 35198 30620 35900 30648
rect 35198 30617 35210 30620
rect 35152 30611 35210 30617
rect 35894 30608 35900 30620
rect 35952 30608 35958 30660
rect 40512 30648 40540 30679
rect 40770 30676 40776 30688
rect 40828 30676 40834 30728
rect 43180 30725 43208 30756
rect 43364 30725 43392 30812
rect 45554 30784 45560 30796
rect 45204 30756 45560 30784
rect 43165 30719 43223 30725
rect 43165 30685 43177 30719
rect 43211 30685 43223 30719
rect 43165 30679 43223 30685
rect 43257 30719 43315 30725
rect 43257 30685 43269 30719
rect 43303 30685 43315 30719
rect 43257 30679 43315 30685
rect 43349 30719 43407 30725
rect 43349 30685 43361 30719
rect 43395 30685 43407 30719
rect 43530 30716 43536 30728
rect 43491 30688 43536 30716
rect 43349 30679 43407 30685
rect 41138 30648 41144 30660
rect 40512 30620 41144 30648
rect 41138 30608 41144 30620
rect 41196 30608 41202 30660
rect 43272 30592 43300 30679
rect 43530 30676 43536 30688
rect 43588 30676 43594 30728
rect 45204 30725 45232 30756
rect 45554 30744 45560 30756
rect 45612 30744 45618 30796
rect 45370 30725 45376 30728
rect 45189 30719 45247 30725
rect 45189 30685 45201 30719
rect 45235 30685 45247 30719
rect 45189 30679 45247 30685
rect 45337 30719 45376 30725
rect 45337 30685 45349 30719
rect 45337 30679 45376 30685
rect 45370 30676 45376 30679
rect 45428 30676 45434 30728
rect 45654 30719 45712 30725
rect 45654 30685 45666 30719
rect 45700 30716 45712 30719
rect 45700 30688 45784 30716
rect 45700 30685 45712 30688
rect 45654 30679 45712 30685
rect 45465 30651 45523 30657
rect 45465 30617 45477 30651
rect 45511 30617 45523 30651
rect 45465 30611 45523 30617
rect 45557 30651 45615 30657
rect 45557 30617 45569 30651
rect 45603 30617 45615 30651
rect 45756 30648 45784 30688
rect 45830 30676 45836 30728
rect 45888 30716 45894 30728
rect 46293 30719 46351 30725
rect 46293 30716 46305 30719
rect 45888 30688 46305 30716
rect 45888 30676 45894 30688
rect 46293 30685 46305 30688
rect 46339 30685 46351 30719
rect 46293 30679 46351 30685
rect 46385 30651 46443 30657
rect 46385 30648 46397 30651
rect 45756 30620 46397 30648
rect 45557 30611 45615 30617
rect 46385 30617 46397 30620
rect 46431 30617 46443 30651
rect 46385 30611 46443 30617
rect 26329 30583 26387 30589
rect 26329 30549 26341 30583
rect 26375 30580 26387 30583
rect 26602 30580 26608 30592
rect 26375 30552 26608 30580
rect 26375 30549 26387 30552
rect 26329 30543 26387 30549
rect 26602 30540 26608 30552
rect 26660 30540 26666 30592
rect 31573 30583 31631 30589
rect 31573 30549 31585 30583
rect 31619 30580 31631 30583
rect 31662 30580 31668 30592
rect 31619 30552 31668 30580
rect 31619 30549 31631 30552
rect 31573 30543 31631 30549
rect 31662 30540 31668 30552
rect 31720 30540 31726 30592
rect 36170 30540 36176 30592
rect 36228 30580 36234 30592
rect 36265 30583 36323 30589
rect 36265 30580 36277 30583
rect 36228 30552 36277 30580
rect 36228 30540 36234 30552
rect 36265 30549 36277 30552
rect 36311 30549 36323 30583
rect 36265 30543 36323 30549
rect 40034 30540 40040 30592
rect 40092 30580 40098 30592
rect 40681 30583 40739 30589
rect 40681 30580 40693 30583
rect 40092 30552 40693 30580
rect 40092 30540 40098 30552
rect 40681 30549 40693 30552
rect 40727 30549 40739 30583
rect 42886 30580 42892 30592
rect 42847 30552 42892 30580
rect 40681 30543 40739 30549
rect 42886 30540 42892 30552
rect 42944 30540 42950 30592
rect 43254 30540 43260 30592
rect 43312 30540 43318 30592
rect 45186 30540 45192 30592
rect 45244 30580 45250 30592
rect 45480 30580 45508 30611
rect 45244 30552 45508 30580
rect 45572 30580 45600 30611
rect 46014 30580 46020 30592
rect 45572 30552 46020 30580
rect 45244 30540 45250 30552
rect 46014 30540 46020 30552
rect 46072 30540 46078 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 23474 30336 23480 30388
rect 23532 30376 23538 30388
rect 25409 30379 25467 30385
rect 25409 30376 25421 30379
rect 23532 30348 25421 30376
rect 23532 30336 23538 30348
rect 25409 30345 25421 30348
rect 25455 30345 25467 30379
rect 25409 30339 25467 30345
rect 26050 30336 26056 30388
rect 26108 30376 26114 30388
rect 30006 30376 30012 30388
rect 26108 30348 30012 30376
rect 26108 30336 26114 30348
rect 30006 30336 30012 30348
rect 30064 30336 30070 30388
rect 33134 30376 33140 30388
rect 33095 30348 33140 30376
rect 33134 30336 33140 30348
rect 33192 30336 33198 30388
rect 40129 30379 40187 30385
rect 40129 30345 40141 30379
rect 40175 30376 40187 30379
rect 40770 30376 40776 30388
rect 40175 30348 40776 30376
rect 40175 30345 40187 30348
rect 40129 30339 40187 30345
rect 40770 30336 40776 30348
rect 40828 30336 40834 30388
rect 41138 30376 41144 30388
rect 41099 30348 41144 30376
rect 41138 30336 41144 30348
rect 41196 30336 41202 30388
rect 42812 30348 43392 30376
rect 23290 30268 23296 30320
rect 23348 30308 23354 30320
rect 26068 30308 26096 30336
rect 23348 30280 26096 30308
rect 23348 30268 23354 30280
rect 31386 30268 31392 30320
rect 31444 30308 31450 30320
rect 36170 30308 36176 30320
rect 31444 30280 32536 30308
rect 31444 30268 31450 30280
rect 23382 30200 23388 30252
rect 23440 30240 23446 30252
rect 24285 30243 24343 30249
rect 24285 30240 24297 30243
rect 23440 30212 24297 30240
rect 23440 30200 23446 30212
rect 24285 30209 24297 30212
rect 24331 30209 24343 30243
rect 31662 30240 31668 30252
rect 31623 30212 31668 30240
rect 24285 30203 24343 30209
rect 31662 30200 31668 30212
rect 31720 30200 31726 30252
rect 32122 30200 32128 30252
rect 32180 30240 32186 30252
rect 32306 30240 32312 30252
rect 32180 30212 32312 30240
rect 32180 30200 32186 30212
rect 32306 30200 32312 30212
rect 32364 30200 32370 30252
rect 32508 30249 32536 30280
rect 35360 30280 36176 30308
rect 35360 30249 35388 30280
rect 36170 30268 36176 30280
rect 36228 30268 36234 30320
rect 39117 30311 39175 30317
rect 39117 30277 39129 30311
rect 39163 30277 39175 30311
rect 39117 30271 39175 30277
rect 39853 30311 39911 30317
rect 39853 30277 39865 30311
rect 39899 30308 39911 30311
rect 40494 30308 40500 30320
rect 39899 30280 40500 30308
rect 39899 30277 39911 30280
rect 39853 30271 39911 30277
rect 32493 30243 32551 30249
rect 32493 30209 32505 30243
rect 32539 30209 32551 30243
rect 32493 30203 32551 30209
rect 32677 30243 32735 30249
rect 32677 30209 32689 30243
rect 32723 30240 32735 30243
rect 33321 30243 33379 30249
rect 33321 30240 33333 30243
rect 32723 30212 33333 30240
rect 32723 30209 32735 30212
rect 32677 30203 32735 30209
rect 33321 30209 33333 30212
rect 33367 30209 33379 30243
rect 33321 30203 33379 30209
rect 35345 30243 35403 30249
rect 35345 30209 35357 30243
rect 35391 30209 35403 30243
rect 35345 30203 35403 30209
rect 35434 30200 35440 30252
rect 35492 30240 35498 30252
rect 35529 30243 35587 30249
rect 35529 30240 35541 30243
rect 35492 30212 35541 30240
rect 35492 30200 35498 30212
rect 35529 30209 35541 30212
rect 35575 30209 35587 30243
rect 38838 30240 38844 30252
rect 38799 30212 38844 30240
rect 35529 30203 35587 30209
rect 38838 30200 38844 30212
rect 38896 30200 38902 30252
rect 39132 30240 39160 30271
rect 40494 30268 40500 30280
rect 40552 30268 40558 30320
rect 40865 30311 40923 30317
rect 40865 30277 40877 30311
rect 40911 30308 40923 30311
rect 41322 30308 41328 30320
rect 40911 30280 41328 30308
rect 40911 30277 40923 30280
rect 40865 30271 40923 30277
rect 41322 30268 41328 30280
rect 41380 30268 41386 30320
rect 39577 30243 39635 30249
rect 39577 30240 39589 30243
rect 39132 30212 39589 30240
rect 39577 30209 39589 30212
rect 39623 30209 39635 30243
rect 39758 30240 39764 30252
rect 39719 30212 39764 30240
rect 39577 30203 39635 30209
rect 39758 30200 39764 30212
rect 39816 30200 39822 30252
rect 39945 30243 40003 30249
rect 39945 30209 39957 30243
rect 39991 30240 40003 30243
rect 40218 30240 40224 30252
rect 39991 30212 40224 30240
rect 39991 30209 40003 30212
rect 39945 30203 40003 30209
rect 40218 30200 40224 30212
rect 40276 30200 40282 30252
rect 40586 30240 40592 30252
rect 40547 30212 40592 30240
rect 40586 30200 40592 30212
rect 40644 30200 40650 30252
rect 40770 30240 40776 30252
rect 40731 30212 40776 30240
rect 40770 30200 40776 30212
rect 40828 30200 40834 30252
rect 40957 30243 41015 30249
rect 40957 30209 40969 30243
rect 41003 30240 41015 30243
rect 41966 30240 41972 30252
rect 41003 30212 41972 30240
rect 41003 30209 41015 30212
rect 40957 30203 41015 30209
rect 41966 30200 41972 30212
rect 42024 30200 42030 30252
rect 24029 30175 24087 30181
rect 24029 30141 24041 30175
rect 24075 30141 24087 30175
rect 24029 30135 24087 30141
rect 39117 30175 39175 30181
rect 39117 30141 39129 30175
rect 39163 30172 39175 30175
rect 42812 30172 42840 30348
rect 42886 30268 42892 30320
rect 42944 30308 42950 30320
rect 43226 30311 43284 30317
rect 43226 30308 43238 30311
rect 42944 30280 43238 30308
rect 42944 30268 42950 30280
rect 43226 30277 43238 30280
rect 43272 30277 43284 30311
rect 43364 30308 43392 30348
rect 43364 30280 45508 30308
rect 43226 30271 43284 30277
rect 43070 30200 43076 30252
rect 43128 30240 43134 30252
rect 44821 30243 44879 30249
rect 44821 30240 44833 30243
rect 43128 30212 44833 30240
rect 43128 30200 43134 30212
rect 44821 30209 44833 30212
rect 44867 30209 44879 30243
rect 45002 30240 45008 30252
rect 44963 30212 45008 30240
rect 44821 30203 44879 30209
rect 45002 30200 45008 30212
rect 45060 30200 45066 30252
rect 45370 30240 45376 30252
rect 45331 30212 45376 30240
rect 45370 30200 45376 30212
rect 45428 30200 45434 30252
rect 39163 30144 42840 30172
rect 39163 30141 39175 30144
rect 39117 30135 39175 30141
rect 24044 30036 24072 30135
rect 42886 30132 42892 30184
rect 42944 30172 42950 30184
rect 42981 30175 43039 30181
rect 42981 30172 42993 30175
rect 42944 30144 42993 30172
rect 42944 30132 42950 30144
rect 42981 30141 42993 30144
rect 43027 30141 43039 30175
rect 45094 30172 45100 30184
rect 45055 30144 45100 30172
rect 42981 30135 43039 30141
rect 45094 30132 45100 30144
rect 45152 30132 45158 30184
rect 45186 30132 45192 30184
rect 45244 30172 45250 30184
rect 45480 30172 45508 30280
rect 45830 30200 45836 30252
rect 45888 30240 45894 30252
rect 46017 30243 46075 30249
rect 46017 30240 46029 30243
rect 45888 30212 46029 30240
rect 45888 30200 45894 30212
rect 46017 30209 46029 30212
rect 46063 30209 46075 30243
rect 46017 30203 46075 30209
rect 47486 30200 47492 30252
rect 47544 30240 47550 30252
rect 47670 30240 47676 30252
rect 47544 30212 47676 30240
rect 47544 30200 47550 30212
rect 47670 30200 47676 30212
rect 47728 30240 47734 30252
rect 47765 30243 47823 30249
rect 47765 30240 47777 30243
rect 47728 30212 47777 30240
rect 47728 30200 47734 30212
rect 47765 30209 47777 30212
rect 47811 30209 47823 30243
rect 47765 30203 47823 30209
rect 46198 30172 46204 30184
rect 45244 30144 45289 30172
rect 45480 30144 46204 30172
rect 45244 30132 45250 30144
rect 46198 30132 46204 30144
rect 46256 30172 46262 30184
rect 46477 30175 46535 30181
rect 46477 30172 46489 30175
rect 46256 30144 46489 30172
rect 46256 30132 46262 30144
rect 46477 30141 46489 30144
rect 46523 30141 46535 30175
rect 46477 30135 46535 30141
rect 44082 30064 44088 30116
rect 44140 30104 44146 30116
rect 44361 30107 44419 30113
rect 44361 30104 44373 30107
rect 44140 30076 44373 30104
rect 44140 30064 44146 30076
rect 44361 30073 44373 30076
rect 44407 30073 44419 30107
rect 44361 30067 44419 30073
rect 24394 30036 24400 30048
rect 24044 30008 24400 30036
rect 24394 29996 24400 30008
rect 24452 29996 24458 30048
rect 31481 30039 31539 30045
rect 31481 30005 31493 30039
rect 31527 30036 31539 30039
rect 31570 30036 31576 30048
rect 31527 30008 31576 30036
rect 31527 30005 31539 30008
rect 31481 29999 31539 30005
rect 31570 29996 31576 30008
rect 31628 29996 31634 30048
rect 35342 30036 35348 30048
rect 35303 30008 35348 30036
rect 35342 29996 35348 30008
rect 35400 29996 35406 30048
rect 38930 30036 38936 30048
rect 38891 30008 38936 30036
rect 38930 29996 38936 30008
rect 38988 29996 38994 30048
rect 43622 29996 43628 30048
rect 43680 30036 43686 30048
rect 44100 30036 44128 30064
rect 45554 30036 45560 30048
rect 43680 30008 44128 30036
rect 45515 30008 45560 30036
rect 43680 29996 43686 30008
rect 45554 29996 45560 30008
rect 45612 29996 45618 30048
rect 46014 29996 46020 30048
rect 46072 30036 46078 30048
rect 46109 30039 46167 30045
rect 46109 30036 46121 30039
rect 46072 30008 46121 30036
rect 46072 29996 46078 30008
rect 46109 30005 46121 30008
rect 46155 30005 46167 30039
rect 47210 30036 47216 30048
rect 47171 30008 47216 30036
rect 46109 29999 46167 30005
rect 47210 29996 47216 30008
rect 47268 29996 47274 30048
rect 47854 30036 47860 30048
rect 47815 30008 47860 30036
rect 47854 29996 47860 30008
rect 47912 29996 47918 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 23382 29832 23388 29844
rect 23343 29804 23388 29832
rect 23382 29792 23388 29804
rect 23440 29792 23446 29844
rect 27430 29792 27436 29844
rect 27488 29832 27494 29844
rect 28629 29835 28687 29841
rect 28629 29832 28641 29835
rect 27488 29804 28641 29832
rect 27488 29792 27494 29804
rect 28629 29801 28641 29804
rect 28675 29801 28687 29835
rect 28629 29795 28687 29801
rect 32306 29792 32312 29844
rect 32364 29832 32370 29844
rect 32677 29835 32735 29841
rect 32677 29832 32689 29835
rect 32364 29804 32689 29832
rect 32364 29792 32370 29804
rect 32677 29801 32689 29804
rect 32723 29801 32735 29835
rect 32677 29795 32735 29801
rect 39025 29835 39083 29841
rect 39025 29801 39037 29835
rect 39071 29832 39083 29835
rect 39758 29832 39764 29844
rect 39071 29804 39764 29832
rect 39071 29801 39083 29804
rect 39025 29795 39083 29801
rect 39758 29792 39764 29804
rect 39816 29792 39822 29844
rect 40034 29832 40040 29844
rect 39995 29804 40040 29832
rect 40034 29792 40040 29804
rect 40092 29792 40098 29844
rect 40497 29835 40555 29841
rect 40497 29801 40509 29835
rect 40543 29832 40555 29835
rect 40770 29832 40776 29844
rect 40543 29804 40776 29832
rect 40543 29801 40555 29804
rect 40497 29795 40555 29801
rect 40770 29792 40776 29804
rect 40828 29792 40834 29844
rect 45186 29792 45192 29844
rect 45244 29832 45250 29844
rect 45741 29835 45799 29841
rect 45741 29832 45753 29835
rect 45244 29804 45753 29832
rect 45244 29792 45250 29804
rect 45741 29801 45753 29804
rect 45787 29801 45799 29835
rect 45741 29795 45799 29801
rect 22833 29767 22891 29773
rect 22833 29733 22845 29767
rect 22879 29764 22891 29767
rect 24762 29764 24768 29776
rect 22879 29736 24768 29764
rect 22879 29733 22891 29736
rect 22833 29727 22891 29733
rect 23676 29696 23704 29736
rect 24762 29724 24768 29736
rect 24820 29724 24826 29776
rect 35434 29764 35440 29776
rect 35176 29736 35440 29764
rect 23676 29668 23796 29696
rect 22649 29631 22707 29637
rect 22649 29597 22661 29631
rect 22695 29628 22707 29631
rect 23290 29628 23296 29640
rect 22695 29600 23296 29628
rect 22695 29597 22707 29600
rect 22649 29591 22707 29597
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 23566 29588 23572 29640
rect 23624 29638 23630 29640
rect 23624 29637 23704 29638
rect 23768 29637 23796 29668
rect 24394 29656 24400 29708
rect 24452 29696 24458 29708
rect 35176 29705 35204 29736
rect 35434 29724 35440 29736
rect 35492 29724 35498 29776
rect 27249 29699 27307 29705
rect 27249 29696 27261 29699
rect 24452 29668 27261 29696
rect 24452 29656 24458 29668
rect 27249 29665 27261 29668
rect 27295 29665 27307 29699
rect 27249 29659 27307 29665
rect 35161 29699 35219 29705
rect 35161 29665 35173 29699
rect 35207 29665 35219 29699
rect 35161 29659 35219 29665
rect 35253 29699 35311 29705
rect 35253 29665 35265 29699
rect 35299 29696 35311 29699
rect 35299 29668 36216 29696
rect 35299 29665 35311 29668
rect 35253 29659 35311 29665
rect 23624 29631 23719 29637
rect 23624 29610 23673 29631
rect 23624 29588 23630 29610
rect 23661 29597 23673 29610
rect 23707 29597 23719 29631
rect 23661 29591 23719 29597
rect 23750 29631 23808 29637
rect 23750 29597 23762 29631
rect 23796 29597 23808 29631
rect 23750 29591 23808 29597
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29597 23903 29631
rect 23845 29591 23903 29597
rect 23860 29492 23888 29591
rect 24026 29588 24032 29640
rect 24084 29628 24090 29640
rect 26329 29631 26387 29637
rect 24084 29600 24129 29628
rect 24084 29588 24090 29600
rect 26329 29597 26341 29631
rect 26375 29597 26387 29631
rect 26602 29628 26608 29640
rect 26563 29600 26608 29628
rect 26329 29591 26387 29597
rect 26344 29560 26372 29591
rect 26602 29588 26608 29600
rect 26660 29588 26666 29640
rect 27264 29628 27292 29659
rect 28718 29628 28724 29640
rect 27264 29600 28724 29628
rect 28718 29588 28724 29600
rect 28776 29588 28782 29640
rect 31570 29637 31576 29640
rect 31297 29631 31355 29637
rect 31297 29597 31309 29631
rect 31343 29597 31355 29631
rect 31564 29628 31576 29637
rect 31531 29600 31576 29628
rect 31297 29591 31355 29597
rect 31564 29591 31576 29600
rect 26418 29560 26424 29572
rect 26331 29532 26424 29560
rect 26418 29520 26424 29532
rect 26476 29560 26482 29572
rect 26476 29532 26648 29560
rect 26476 29520 26482 29532
rect 23934 29492 23940 29504
rect 23860 29464 23940 29492
rect 23934 29452 23940 29464
rect 23992 29452 23998 29504
rect 24578 29452 24584 29504
rect 24636 29492 24642 29504
rect 26145 29495 26203 29501
rect 26145 29492 26157 29495
rect 24636 29464 26157 29492
rect 24636 29452 24642 29464
rect 26145 29461 26157 29464
rect 26191 29461 26203 29495
rect 26510 29492 26516 29504
rect 26471 29464 26516 29492
rect 26145 29455 26203 29461
rect 26510 29452 26516 29464
rect 26568 29452 26574 29504
rect 26620 29492 26648 29532
rect 27154 29520 27160 29572
rect 27212 29560 27218 29572
rect 27494 29563 27552 29569
rect 27494 29560 27506 29563
rect 27212 29532 27506 29560
rect 27212 29520 27218 29532
rect 27494 29529 27506 29532
rect 27540 29529 27552 29563
rect 27494 29523 27552 29529
rect 27890 29492 27896 29504
rect 26620 29464 27896 29492
rect 27890 29452 27896 29464
rect 27948 29452 27954 29504
rect 31312 29492 31340 29591
rect 31570 29588 31576 29591
rect 31628 29588 31634 29640
rect 34238 29588 34244 29640
rect 34296 29628 34302 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34296 29600 34897 29628
rect 34296 29588 34302 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 35176 29628 35204 29659
rect 36188 29640 36216 29668
rect 38838 29656 38844 29708
rect 38896 29696 38902 29708
rect 38896 29668 39160 29696
rect 38896 29656 38902 29668
rect 35989 29631 36047 29637
rect 35989 29628 36001 29631
rect 35176 29600 36001 29628
rect 34885 29591 34943 29597
rect 35989 29597 36001 29600
rect 36035 29597 36047 29631
rect 36170 29628 36176 29640
rect 36131 29600 36176 29628
rect 35989 29591 36047 29597
rect 36170 29588 36176 29600
rect 36228 29588 36234 29640
rect 38930 29628 38936 29640
rect 38891 29600 38936 29628
rect 38930 29588 38936 29600
rect 38988 29588 38994 29640
rect 39132 29637 39160 29668
rect 41322 29656 41328 29708
rect 41380 29696 41386 29708
rect 42981 29699 43039 29705
rect 41380 29668 42840 29696
rect 41380 29656 41386 29668
rect 39117 29631 39175 29637
rect 39117 29597 39129 29631
rect 39163 29597 39175 29631
rect 40218 29628 40224 29640
rect 40179 29600 40224 29628
rect 39117 29591 39175 29597
rect 40218 29588 40224 29600
rect 40276 29588 40282 29640
rect 40313 29631 40371 29637
rect 40313 29597 40325 29631
rect 40359 29628 40371 29631
rect 40494 29628 40500 29640
rect 40359 29600 40500 29628
rect 40359 29597 40371 29600
rect 40313 29591 40371 29597
rect 40494 29588 40500 29600
rect 40552 29588 40558 29640
rect 40586 29588 40592 29640
rect 40644 29628 40650 29640
rect 40644 29600 40689 29628
rect 40644 29588 40650 29600
rect 41966 29588 41972 29640
rect 42024 29628 42030 29640
rect 42812 29637 42840 29668
rect 42981 29665 42993 29699
rect 43027 29696 43039 29699
rect 46477 29699 46535 29705
rect 43027 29668 43760 29696
rect 43027 29665 43039 29668
rect 42981 29659 43039 29665
rect 43732 29640 43760 29668
rect 46477 29665 46489 29699
rect 46523 29696 46535 29699
rect 47210 29696 47216 29708
rect 46523 29668 47216 29696
rect 46523 29665 46535 29668
rect 46477 29659 46535 29665
rect 47210 29656 47216 29668
rect 47268 29656 47274 29708
rect 42705 29631 42763 29637
rect 42705 29628 42717 29631
rect 42024 29600 42717 29628
rect 42024 29588 42030 29600
rect 42705 29597 42717 29600
rect 42751 29597 42763 29631
rect 42705 29591 42763 29597
rect 42797 29631 42855 29637
rect 42797 29597 42809 29631
rect 42843 29597 42855 29631
rect 42797 29591 42855 29597
rect 43073 29631 43131 29637
rect 43073 29597 43085 29631
rect 43119 29628 43131 29631
rect 43533 29631 43591 29637
rect 43533 29628 43545 29631
rect 43119 29600 43545 29628
rect 43119 29597 43131 29600
rect 43073 29591 43131 29597
rect 43533 29597 43545 29600
rect 43579 29628 43591 29631
rect 43622 29628 43628 29640
rect 43579 29600 43628 29628
rect 43579 29597 43591 29600
rect 43533 29591 43591 29597
rect 43622 29588 43628 29600
rect 43680 29588 43686 29640
rect 43714 29588 43720 29640
rect 43772 29628 43778 29640
rect 43901 29631 43959 29637
rect 43772 29600 43865 29628
rect 43772 29588 43778 29600
rect 43901 29597 43913 29631
rect 43947 29628 43959 29631
rect 43990 29628 43996 29640
rect 43947 29600 43996 29628
rect 43947 29597 43959 29600
rect 43901 29591 43959 29597
rect 43990 29588 43996 29600
rect 44048 29628 44054 29640
rect 45002 29628 45008 29640
rect 44048 29600 45008 29628
rect 44048 29588 44054 29600
rect 45002 29588 45008 29600
rect 45060 29588 45066 29640
rect 45649 29631 45707 29637
rect 45649 29597 45661 29631
rect 45695 29628 45707 29631
rect 45738 29628 45744 29640
rect 45695 29600 45744 29628
rect 45695 29597 45707 29600
rect 45649 29591 45707 29597
rect 45738 29588 45744 29600
rect 45796 29588 45802 29640
rect 34606 29520 34612 29572
rect 34664 29560 34670 29572
rect 35370 29563 35428 29569
rect 35370 29560 35382 29563
rect 34664 29532 35382 29560
rect 34664 29520 34670 29532
rect 35370 29529 35382 29532
rect 35416 29560 35428 29563
rect 35618 29560 35624 29572
rect 35416 29532 35624 29560
rect 35416 29529 35428 29532
rect 35370 29523 35428 29529
rect 35618 29520 35624 29532
rect 35676 29520 35682 29572
rect 43809 29563 43867 29569
rect 43809 29529 43821 29563
rect 43855 29560 43867 29563
rect 45094 29560 45100 29572
rect 43855 29532 45100 29560
rect 43855 29529 43867 29532
rect 43809 29523 43867 29529
rect 45094 29520 45100 29532
rect 45152 29520 45158 29572
rect 46661 29563 46719 29569
rect 46661 29529 46673 29563
rect 46707 29560 46719 29563
rect 47854 29560 47860 29572
rect 46707 29532 47860 29560
rect 46707 29529 46719 29532
rect 46661 29523 46719 29529
rect 47854 29520 47860 29532
rect 47912 29520 47918 29572
rect 48314 29560 48320 29572
rect 48275 29532 48320 29560
rect 48314 29520 48320 29532
rect 48372 29520 48378 29572
rect 31754 29492 31760 29504
rect 31312 29464 31760 29492
rect 31754 29452 31760 29464
rect 31812 29492 31818 29504
rect 32214 29492 32220 29504
rect 31812 29464 32220 29492
rect 31812 29452 31818 29464
rect 32214 29452 32220 29464
rect 32272 29452 32278 29504
rect 35529 29495 35587 29501
rect 35529 29461 35541 29495
rect 35575 29492 35587 29495
rect 35894 29492 35900 29504
rect 35575 29464 35900 29492
rect 35575 29461 35587 29464
rect 35529 29455 35587 29461
rect 35894 29452 35900 29464
rect 35952 29452 35958 29504
rect 36354 29492 36360 29504
rect 36315 29464 36360 29492
rect 36354 29452 36360 29464
rect 36412 29452 36418 29504
rect 42521 29495 42579 29501
rect 42521 29461 42533 29495
rect 42567 29492 42579 29495
rect 43254 29492 43260 29504
rect 42567 29464 43260 29492
rect 42567 29461 42579 29464
rect 42521 29455 42579 29461
rect 43254 29452 43260 29464
rect 43312 29452 43318 29504
rect 44082 29492 44088 29504
rect 44043 29464 44088 29492
rect 44082 29452 44088 29464
rect 44140 29452 44146 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 23290 29288 23296 29300
rect 23251 29260 23296 29288
rect 23290 29248 23296 29260
rect 23348 29248 23354 29300
rect 23934 29288 23940 29300
rect 23895 29260 23940 29288
rect 23934 29248 23940 29260
rect 23992 29248 23998 29300
rect 24026 29248 24032 29300
rect 24084 29288 24090 29300
rect 27154 29288 27160 29300
rect 24084 29260 27016 29288
rect 27115 29260 27160 29288
rect 24084 29248 24090 29260
rect 24670 29220 24676 29232
rect 24412 29192 24676 29220
rect 24412 29161 24440 29192
rect 24670 29180 24676 29192
rect 24728 29180 24734 29232
rect 26988 29220 27016 29260
rect 27154 29248 27160 29260
rect 27212 29248 27218 29300
rect 27816 29260 35664 29288
rect 27816 29220 27844 29260
rect 29362 29220 29368 29232
rect 26988 29192 27844 29220
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29121 24455 29155
rect 24578 29152 24584 29164
rect 24539 29124 24584 29152
rect 24397 29115 24455 29121
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 26418 29152 26424 29164
rect 26379 29124 26424 29152
rect 26418 29112 26424 29124
rect 26476 29112 26482 29164
rect 26602 29152 26608 29164
rect 26563 29124 26608 29152
rect 26602 29112 26608 29124
rect 26660 29112 26666 29164
rect 27430 29152 27436 29164
rect 27391 29124 27436 29152
rect 27430 29112 27436 29124
rect 27488 29112 27494 29164
rect 27525 29155 27583 29161
rect 27525 29121 27537 29155
rect 27571 29121 27583 29155
rect 27525 29115 27583 29121
rect 23658 29084 23664 29096
rect 23619 29056 23664 29084
rect 23658 29044 23664 29056
rect 23716 29044 23722 29096
rect 23753 29087 23811 29093
rect 23753 29053 23765 29087
rect 23799 29084 23811 29087
rect 23799 29056 24532 29084
rect 23799 29053 23811 29056
rect 23753 29047 23811 29053
rect 24504 28960 24532 29056
rect 24762 29044 24768 29096
rect 24820 29084 24826 29096
rect 27540 29084 27568 29115
rect 27614 29112 27620 29164
rect 27672 29152 27678 29164
rect 27816 29161 27844 29192
rect 28736 29192 29368 29220
rect 28736 29164 28764 29192
rect 29362 29180 29368 29192
rect 29420 29220 29426 29232
rect 29822 29220 29828 29232
rect 29420 29192 29828 29220
rect 29420 29180 29426 29192
rect 29822 29180 29828 29192
rect 29880 29180 29886 29232
rect 33410 29180 33416 29232
rect 33468 29220 33474 29232
rect 34238 29220 34244 29232
rect 33468 29192 34244 29220
rect 33468 29180 33474 29192
rect 34238 29180 34244 29192
rect 34296 29220 34302 29232
rect 35636 29220 35664 29260
rect 35710 29248 35716 29300
rect 35768 29288 35774 29300
rect 40129 29291 40187 29297
rect 35768 29260 36216 29288
rect 35768 29248 35774 29260
rect 36188 29229 36216 29260
rect 40129 29257 40141 29291
rect 40175 29288 40187 29291
rect 40218 29288 40224 29300
rect 40175 29260 40224 29288
rect 40175 29257 40187 29260
rect 40129 29251 40187 29257
rect 40218 29248 40224 29260
rect 40276 29248 40282 29300
rect 40770 29288 40776 29300
rect 40731 29260 40776 29288
rect 40770 29248 40776 29260
rect 40828 29248 40834 29300
rect 41966 29288 41972 29300
rect 41927 29260 41972 29288
rect 41966 29248 41972 29260
rect 42024 29248 42030 29300
rect 42889 29291 42947 29297
rect 42889 29257 42901 29291
rect 42935 29288 42947 29291
rect 43070 29288 43076 29300
rect 42935 29260 43076 29288
rect 42935 29257 42947 29260
rect 42889 29251 42947 29257
rect 43070 29248 43076 29260
rect 43128 29248 43134 29300
rect 43254 29288 43260 29300
rect 43215 29260 43260 29288
rect 43254 29248 43260 29260
rect 43312 29248 43318 29300
rect 43714 29248 43720 29300
rect 43772 29288 43778 29300
rect 43901 29291 43959 29297
rect 43901 29288 43913 29291
rect 43772 29260 43913 29288
rect 43772 29248 43778 29260
rect 43901 29257 43913 29260
rect 43947 29257 43959 29291
rect 43901 29251 43959 29257
rect 36173 29223 36231 29229
rect 34296 29192 35572 29220
rect 35636 29192 36124 29220
rect 34296 29180 34302 29192
rect 27801 29155 27859 29161
rect 27672 29124 27717 29152
rect 27672 29112 27678 29124
rect 27801 29121 27813 29155
rect 27847 29121 27859 29155
rect 28718 29152 28724 29164
rect 28679 29124 28724 29152
rect 27801 29115 27859 29121
rect 28718 29112 28724 29124
rect 28776 29112 28782 29164
rect 28988 29155 29046 29161
rect 28988 29121 29000 29155
rect 29034 29152 29046 29155
rect 30561 29155 30619 29161
rect 30561 29152 30573 29155
rect 29034 29124 30573 29152
rect 29034 29121 29046 29124
rect 28988 29115 29046 29121
rect 30561 29121 30573 29124
rect 30607 29121 30619 29155
rect 30742 29152 30748 29164
rect 30703 29124 30748 29152
rect 30561 29115 30619 29121
rect 30742 29112 30748 29124
rect 30800 29112 30806 29164
rect 35342 29152 35348 29164
rect 35303 29124 35348 29152
rect 35342 29112 35348 29124
rect 35400 29112 35406 29164
rect 35437 29155 35495 29161
rect 35437 29121 35449 29155
rect 35483 29121 35495 29155
rect 35437 29115 35495 29121
rect 24820 29056 27660 29084
rect 24820 29044 24826 29056
rect 24486 28948 24492 28960
rect 24447 28920 24492 28948
rect 24486 28908 24492 28920
rect 24544 28908 24550 28960
rect 26421 28951 26479 28957
rect 26421 28917 26433 28951
rect 26467 28948 26479 28951
rect 26786 28948 26792 28960
rect 26467 28920 26792 28948
rect 26467 28917 26479 28920
rect 26421 28911 26479 28917
rect 26786 28908 26792 28920
rect 26844 28908 26850 28960
rect 27632 28948 27660 29056
rect 29914 29044 29920 29096
rect 29972 29084 29978 29096
rect 31021 29087 31079 29093
rect 31021 29084 31033 29087
rect 29972 29056 31033 29084
rect 29972 29044 29978 29056
rect 31021 29053 31033 29056
rect 31067 29053 31079 29087
rect 35452 29084 35480 29115
rect 31021 29047 31079 29053
rect 35360 29056 35480 29084
rect 30929 29019 30987 29025
rect 30929 29016 30941 29019
rect 29656 28988 30941 29016
rect 27890 28948 27896 28960
rect 27632 28920 27896 28948
rect 27890 28908 27896 28920
rect 27948 28948 27954 28960
rect 29656 28948 29684 28988
rect 30929 28985 30941 28988
rect 30975 28985 30987 29019
rect 34606 29016 34612 29028
rect 34567 28988 34612 29016
rect 30929 28979 30987 28985
rect 34606 28976 34612 28988
rect 34664 28976 34670 29028
rect 27948 28920 29684 28948
rect 27948 28908 27954 28920
rect 29914 28908 29920 28960
rect 29972 28948 29978 28960
rect 30101 28951 30159 28957
rect 30101 28948 30113 28951
rect 29972 28920 30113 28948
rect 29972 28908 29978 28920
rect 30101 28917 30113 28920
rect 30147 28917 30159 28951
rect 34698 28948 34704 28960
rect 34659 28920 34704 28948
rect 30101 28911 30159 28917
rect 34698 28908 34704 28920
rect 34756 28908 34762 28960
rect 35161 28951 35219 28957
rect 35161 28917 35173 28951
rect 35207 28948 35219 28951
rect 35250 28948 35256 28960
rect 35207 28920 35256 28948
rect 35207 28917 35219 28920
rect 35161 28911 35219 28917
rect 35250 28908 35256 28920
rect 35308 28908 35314 28960
rect 35360 28948 35388 29056
rect 35544 29016 35572 29192
rect 35621 29155 35679 29161
rect 35621 29121 35633 29155
rect 35667 29121 35679 29155
rect 35621 29115 35679 29121
rect 35713 29155 35771 29161
rect 35713 29121 35725 29155
rect 35759 29152 35771 29155
rect 35986 29152 35992 29164
rect 35759 29124 35992 29152
rect 35759 29121 35771 29124
rect 35713 29115 35771 29121
rect 35636 29084 35664 29115
rect 35986 29112 35992 29124
rect 36044 29112 36050 29164
rect 36096 29152 36124 29192
rect 36173 29189 36185 29223
rect 36219 29189 36231 29223
rect 38746 29220 38752 29232
rect 36173 29183 36231 29189
rect 36280 29192 38752 29220
rect 36280 29152 36308 29192
rect 38746 29180 38752 29192
rect 38804 29180 38810 29232
rect 44082 29220 44088 29232
rect 43088 29192 44088 29220
rect 36096 29124 36308 29152
rect 37728 29155 37786 29161
rect 37728 29121 37740 29155
rect 37774 29152 37786 29155
rect 38010 29152 38016 29164
rect 37774 29124 38016 29152
rect 37774 29121 37786 29124
rect 37728 29115 37786 29121
rect 38010 29112 38016 29124
rect 38068 29112 38074 29164
rect 40037 29155 40095 29161
rect 40037 29121 40049 29155
rect 40083 29121 40095 29155
rect 40678 29152 40684 29164
rect 40639 29124 40684 29152
rect 40037 29115 40095 29121
rect 35894 29084 35900 29096
rect 35636 29056 35900 29084
rect 35894 29044 35900 29056
rect 35952 29044 35958 29096
rect 37458 29084 37464 29096
rect 37371 29056 37464 29084
rect 37458 29044 37464 29056
rect 37516 29044 37522 29096
rect 40052 29084 40080 29115
rect 40678 29112 40684 29124
rect 40736 29112 40742 29164
rect 41506 29112 41512 29164
rect 41564 29152 41570 29164
rect 43088 29161 43116 29192
rect 44082 29180 44088 29192
rect 44140 29180 44146 29232
rect 41877 29155 41935 29161
rect 41877 29152 41889 29155
rect 41564 29124 41889 29152
rect 41564 29112 41570 29124
rect 41877 29121 41889 29124
rect 41923 29121 41935 29155
rect 41877 29115 41935 29121
rect 43073 29155 43131 29161
rect 43073 29121 43085 29155
rect 43119 29121 43131 29155
rect 43073 29115 43131 29121
rect 43349 29155 43407 29161
rect 43349 29121 43361 29155
rect 43395 29121 43407 29155
rect 43349 29115 43407 29121
rect 43809 29155 43867 29161
rect 43809 29121 43821 29155
rect 43855 29152 43867 29155
rect 43898 29152 43904 29164
rect 43855 29124 43904 29152
rect 43855 29121 43867 29124
rect 43809 29115 43867 29121
rect 40218 29084 40224 29096
rect 40052 29056 40224 29084
rect 40218 29044 40224 29056
rect 40276 29044 40282 29096
rect 42334 29044 42340 29096
rect 42392 29084 42398 29096
rect 43364 29084 43392 29115
rect 43898 29112 43904 29124
rect 43956 29112 43962 29164
rect 45646 29112 45652 29164
rect 45704 29152 45710 29164
rect 45813 29155 45871 29161
rect 45813 29152 45825 29155
rect 45704 29124 45825 29152
rect 45704 29112 45710 29124
rect 45813 29121 45825 29124
rect 45859 29121 45871 29155
rect 45813 29115 45871 29121
rect 45554 29084 45560 29096
rect 42392 29056 43392 29084
rect 45515 29056 45560 29084
rect 42392 29044 42398 29056
rect 45554 29044 45560 29056
rect 45612 29044 45618 29096
rect 36449 29019 36507 29025
rect 36449 29016 36461 29019
rect 35544 28988 36461 29016
rect 36449 28985 36461 28988
rect 36495 28985 36507 29019
rect 36449 28979 36507 28985
rect 36630 28948 36636 28960
rect 35360 28920 36636 28948
rect 36630 28908 36636 28920
rect 36688 28908 36694 28960
rect 37476 28948 37504 29044
rect 38841 29019 38899 29025
rect 38841 28985 38853 29019
rect 38887 29016 38899 29019
rect 38930 29016 38936 29028
rect 38887 28988 38936 29016
rect 38887 28985 38899 28988
rect 38841 28979 38899 28985
rect 38930 28976 38936 28988
rect 38988 29016 38994 29028
rect 40402 29016 40408 29028
rect 38988 28988 40408 29016
rect 38988 28976 38994 28988
rect 40402 28976 40408 28988
rect 40460 28976 40466 29028
rect 46937 29019 46995 29025
rect 46937 29016 46949 29019
rect 46492 28988 46949 29016
rect 38470 28948 38476 28960
rect 37476 28920 38476 28948
rect 38470 28908 38476 28920
rect 38528 28908 38534 28960
rect 45830 28908 45836 28960
rect 45888 28948 45894 28960
rect 46492 28948 46520 28988
rect 46937 28985 46949 28988
rect 46983 28985 46995 29019
rect 46937 28979 46995 28985
rect 47946 28948 47952 28960
rect 45888 28920 46520 28948
rect 47907 28920 47952 28948
rect 45888 28908 45894 28920
rect 47946 28908 47952 28920
rect 48004 28908 48010 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 23658 28704 23664 28756
rect 23716 28744 23722 28756
rect 24949 28747 25007 28753
rect 24949 28744 24961 28747
rect 23716 28716 24961 28744
rect 23716 28704 23722 28716
rect 24949 28713 24961 28716
rect 24995 28713 25007 28747
rect 24949 28707 25007 28713
rect 26053 28747 26111 28753
rect 26053 28713 26065 28747
rect 26099 28744 26111 28747
rect 26602 28744 26608 28756
rect 26099 28716 26608 28744
rect 26099 28713 26111 28716
rect 26053 28707 26111 28713
rect 26602 28704 26608 28716
rect 26660 28704 26666 28756
rect 27614 28704 27620 28756
rect 27672 28744 27678 28756
rect 27801 28747 27859 28753
rect 27801 28744 27813 28747
rect 27672 28716 27813 28744
rect 27672 28704 27678 28716
rect 27801 28713 27813 28716
rect 27847 28713 27859 28747
rect 27801 28707 27859 28713
rect 29733 28747 29791 28753
rect 29733 28713 29745 28747
rect 29779 28744 29791 28747
rect 30742 28744 30748 28756
rect 29779 28716 30748 28744
rect 29779 28713 29791 28716
rect 29733 28707 29791 28713
rect 30742 28704 30748 28716
rect 30800 28704 30806 28756
rect 35986 28744 35992 28756
rect 35176 28716 35992 28744
rect 26694 28676 26700 28688
rect 23676 28648 26700 28676
rect 23676 28620 23704 28648
rect 26694 28636 26700 28648
rect 26752 28636 26758 28688
rect 27249 28679 27307 28685
rect 27249 28645 27261 28679
rect 27295 28645 27307 28679
rect 27249 28639 27307 28645
rect 23658 28568 23664 28620
rect 23716 28568 23722 28620
rect 24578 28568 24584 28620
rect 24636 28608 24642 28620
rect 26786 28608 26792 28620
rect 24636 28580 24808 28608
rect 26747 28580 26792 28608
rect 24636 28568 24642 28580
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28509 23259 28543
rect 23201 28503 23259 28509
rect 23477 28543 23535 28549
rect 23477 28509 23489 28543
rect 23523 28540 23535 28543
rect 24486 28540 24492 28552
rect 23523 28512 24492 28540
rect 23523 28509 23535 28512
rect 23477 28503 23535 28509
rect 23216 28472 23244 28503
rect 24486 28500 24492 28512
rect 24544 28500 24550 28552
rect 24780 28549 24808 28580
rect 26786 28568 26792 28580
rect 26844 28568 26850 28620
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 26053 28543 26111 28549
rect 26053 28509 26065 28543
rect 26099 28509 26111 28543
rect 26053 28503 26111 28509
rect 26237 28543 26295 28549
rect 26237 28509 26249 28543
rect 26283 28509 26295 28543
rect 26237 28503 26295 28509
rect 24581 28475 24639 28481
rect 23216 28444 23520 28472
rect 22646 28364 22652 28416
rect 22704 28404 22710 28416
rect 23017 28407 23075 28413
rect 23017 28404 23029 28407
rect 22704 28376 23029 28404
rect 22704 28364 22710 28376
rect 23017 28373 23029 28376
rect 23063 28373 23075 28407
rect 23382 28404 23388 28416
rect 23343 28376 23388 28404
rect 23017 28367 23075 28373
rect 23382 28364 23388 28376
rect 23440 28364 23446 28416
rect 23492 28404 23520 28444
rect 24581 28441 24593 28475
rect 24627 28472 24639 28475
rect 24670 28472 24676 28484
rect 24627 28444 24676 28472
rect 24627 28441 24639 28444
rect 24581 28435 24639 28441
rect 24670 28432 24676 28444
rect 24728 28432 24734 28484
rect 24946 28404 24952 28416
rect 23492 28376 24952 28404
rect 24946 28364 24952 28376
rect 25004 28364 25010 28416
rect 26068 28404 26096 28503
rect 26252 28472 26280 28503
rect 26510 28500 26516 28552
rect 26568 28540 26574 28552
rect 26881 28543 26939 28549
rect 26881 28540 26893 28543
rect 26568 28512 26893 28540
rect 26568 28500 26574 28512
rect 26881 28509 26893 28512
rect 26927 28509 26939 28543
rect 27264 28540 27292 28639
rect 27709 28543 27767 28549
rect 27709 28540 27721 28543
rect 27264 28512 27721 28540
rect 26881 28503 26939 28509
rect 27709 28509 27721 28512
rect 27755 28509 27767 28543
rect 27890 28540 27896 28552
rect 27851 28512 27896 28540
rect 27709 28503 27767 28509
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 30006 28540 30012 28552
rect 29967 28512 30012 28540
rect 30006 28500 30012 28512
rect 30064 28500 30070 28552
rect 31205 28543 31263 28549
rect 31205 28509 31217 28543
rect 31251 28540 31263 28543
rect 31754 28540 31760 28552
rect 31251 28512 31760 28540
rect 31251 28509 31263 28512
rect 31205 28503 31263 28509
rect 31754 28500 31760 28512
rect 31812 28500 31818 28552
rect 35176 28549 35204 28716
rect 35986 28704 35992 28716
rect 36044 28744 36050 28756
rect 36906 28744 36912 28756
rect 36044 28716 36912 28744
rect 36044 28704 36050 28716
rect 36906 28704 36912 28716
rect 36964 28704 36970 28756
rect 43990 28704 43996 28756
rect 44048 28744 44054 28756
rect 44085 28747 44143 28753
rect 44085 28744 44097 28747
rect 44048 28716 44097 28744
rect 44048 28704 44054 28716
rect 44085 28713 44097 28716
rect 44131 28713 44143 28747
rect 44085 28707 44143 28713
rect 45557 28747 45615 28753
rect 45557 28713 45569 28747
rect 45603 28744 45615 28747
rect 45646 28744 45652 28756
rect 45603 28716 45652 28744
rect 45603 28713 45615 28716
rect 45557 28707 45615 28713
rect 45646 28704 45652 28716
rect 45704 28704 45710 28756
rect 36354 28676 36360 28688
rect 35544 28648 36360 28676
rect 35434 28608 35440 28620
rect 35268 28580 35440 28608
rect 35161 28543 35219 28549
rect 35161 28509 35173 28543
rect 35207 28509 35219 28543
rect 35161 28503 35219 28509
rect 27430 28472 27436 28484
rect 26252 28444 27436 28472
rect 27430 28432 27436 28444
rect 27488 28432 27494 28484
rect 29733 28475 29791 28481
rect 29733 28441 29745 28475
rect 29779 28472 29791 28475
rect 30650 28472 30656 28484
rect 29779 28444 30656 28472
rect 29779 28441 29791 28444
rect 29733 28435 29791 28441
rect 30650 28432 30656 28444
rect 30708 28432 30714 28484
rect 31472 28475 31530 28481
rect 31472 28441 31484 28475
rect 31518 28472 31530 28475
rect 32950 28472 32956 28484
rect 31518 28444 32956 28472
rect 31518 28441 31530 28444
rect 31472 28435 31530 28441
rect 32950 28432 32956 28444
rect 33008 28432 33014 28484
rect 34698 28432 34704 28484
rect 34756 28472 34762 28484
rect 35268 28472 35296 28580
rect 35434 28568 35440 28580
rect 35492 28568 35498 28620
rect 35544 28617 35572 28648
rect 36354 28636 36360 28648
rect 36412 28636 36418 28688
rect 39206 28636 39212 28688
rect 39264 28676 39270 28688
rect 40037 28679 40095 28685
rect 40037 28676 40049 28679
rect 39264 28648 40049 28676
rect 39264 28636 39270 28648
rect 40037 28645 40049 28648
rect 40083 28645 40095 28679
rect 46842 28676 46848 28688
rect 40037 28639 40095 28645
rect 43364 28648 46848 28676
rect 35529 28611 35587 28617
rect 35529 28577 35541 28611
rect 35575 28577 35587 28611
rect 35986 28608 35992 28620
rect 35529 28571 35587 28577
rect 35728 28580 35992 28608
rect 35345 28543 35403 28549
rect 35345 28509 35357 28543
rect 35391 28540 35403 28543
rect 35618 28540 35624 28552
rect 35391 28512 35624 28540
rect 35391 28509 35403 28512
rect 35345 28503 35403 28509
rect 35618 28500 35624 28512
rect 35676 28500 35682 28552
rect 35728 28549 35756 28580
rect 35986 28568 35992 28580
rect 36044 28608 36050 28620
rect 40126 28608 40132 28620
rect 36044 28580 36676 28608
rect 40039 28580 40132 28608
rect 36044 28568 36050 28580
rect 36648 28552 36676 28580
rect 35713 28543 35771 28549
rect 35713 28509 35725 28543
rect 35759 28509 35771 28543
rect 35713 28503 35771 28509
rect 35894 28500 35900 28552
rect 35952 28540 35958 28552
rect 36541 28543 36599 28549
rect 36541 28540 36553 28543
rect 35952 28512 36553 28540
rect 35952 28500 35958 28512
rect 36541 28509 36553 28512
rect 36587 28509 36599 28543
rect 36541 28503 36599 28509
rect 36630 28500 36636 28552
rect 36688 28540 36694 28552
rect 40052 28549 40080 28580
rect 40126 28568 40132 28580
rect 40184 28608 40190 28620
rect 40678 28608 40684 28620
rect 40184 28580 40684 28608
rect 40184 28568 40190 28580
rect 40678 28568 40684 28580
rect 40736 28568 40742 28620
rect 41138 28568 41144 28620
rect 41196 28608 41202 28620
rect 41785 28611 41843 28617
rect 41785 28608 41797 28611
rect 41196 28580 41797 28608
rect 41196 28568 41202 28580
rect 41785 28577 41797 28580
rect 41831 28608 41843 28611
rect 43364 28608 43392 28648
rect 46842 28636 46848 28648
rect 46900 28636 46906 28688
rect 41831 28580 43392 28608
rect 41831 28577 41843 28580
rect 41785 28571 41843 28577
rect 45830 28568 45836 28620
rect 45888 28608 45894 28620
rect 46017 28611 46075 28617
rect 46017 28608 46029 28611
rect 45888 28580 46029 28608
rect 45888 28568 45894 28580
rect 46017 28577 46029 28580
rect 46063 28577 46075 28611
rect 46017 28571 46075 28577
rect 46477 28611 46535 28617
rect 46477 28577 46489 28611
rect 46523 28608 46535 28611
rect 47946 28608 47952 28620
rect 46523 28580 47952 28608
rect 46523 28577 46535 28580
rect 46477 28571 46535 28577
rect 47946 28568 47952 28580
rect 48004 28568 48010 28620
rect 48222 28608 48228 28620
rect 48183 28580 48228 28608
rect 48222 28568 48228 28580
rect 48280 28568 48286 28620
rect 36725 28543 36783 28549
rect 36725 28540 36737 28543
rect 36688 28512 36737 28540
rect 36688 28500 36694 28512
rect 36725 28509 36737 28512
rect 36771 28509 36783 28543
rect 36725 28503 36783 28509
rect 36817 28543 36875 28549
rect 36817 28509 36829 28543
rect 36863 28509 36875 28543
rect 36817 28503 36875 28509
rect 40037 28543 40095 28549
rect 40037 28509 40049 28543
rect 40083 28509 40095 28543
rect 40218 28540 40224 28552
rect 40179 28512 40224 28540
rect 40037 28503 40095 28509
rect 34756 28444 35296 28472
rect 35636 28472 35664 28500
rect 36832 28472 36860 28503
rect 40218 28500 40224 28512
rect 40276 28500 40282 28552
rect 40313 28543 40371 28549
rect 40313 28509 40325 28543
rect 40359 28540 40371 28543
rect 40402 28540 40408 28552
rect 40359 28512 40408 28540
rect 40359 28509 40371 28512
rect 40313 28503 40371 28509
rect 40402 28500 40408 28512
rect 40460 28500 40466 28552
rect 41506 28540 41512 28552
rect 41467 28512 41512 28540
rect 41506 28500 41512 28512
rect 41564 28500 41570 28552
rect 41598 28500 41604 28552
rect 41656 28540 41662 28552
rect 42245 28543 42303 28549
rect 42245 28540 42257 28543
rect 41656 28512 41701 28540
rect 41800 28512 42257 28540
rect 41656 28500 41662 28512
rect 41800 28481 41828 28512
rect 42245 28509 42257 28512
rect 42291 28509 42303 28543
rect 42426 28540 42432 28552
rect 42387 28512 42432 28540
rect 42245 28503 42303 28509
rect 42426 28500 42432 28512
rect 42484 28500 42490 28552
rect 43806 28500 43812 28552
rect 43864 28540 43870 28552
rect 43993 28543 44051 28549
rect 43993 28540 44005 28543
rect 43864 28512 44005 28540
rect 43864 28500 43870 28512
rect 43993 28509 44005 28512
rect 44039 28509 44051 28543
rect 45738 28540 45744 28552
rect 45699 28512 45744 28540
rect 43993 28503 44051 28509
rect 45738 28500 45744 28512
rect 45796 28500 45802 28552
rect 45922 28540 45928 28552
rect 45883 28512 45928 28540
rect 45922 28500 45928 28512
rect 45980 28500 45986 28552
rect 35636 28444 36860 28472
rect 41785 28475 41843 28481
rect 34756 28432 34762 28444
rect 41785 28441 41797 28475
rect 41831 28441 41843 28475
rect 41785 28435 41843 28441
rect 46661 28475 46719 28481
rect 46661 28441 46673 28475
rect 46707 28472 46719 28475
rect 47854 28472 47860 28484
rect 46707 28444 47860 28472
rect 46707 28441 46719 28444
rect 46661 28435 46719 28441
rect 47854 28432 47860 28444
rect 47912 28432 47918 28484
rect 26602 28404 26608 28416
rect 26068 28376 26608 28404
rect 26602 28364 26608 28376
rect 26660 28364 26666 28416
rect 29914 28404 29920 28416
rect 29875 28376 29920 28404
rect 29914 28364 29920 28376
rect 29972 28364 29978 28416
rect 32306 28364 32312 28416
rect 32364 28404 32370 28416
rect 32585 28407 32643 28413
rect 32585 28404 32597 28407
rect 32364 28376 32597 28404
rect 32364 28364 32370 28376
rect 32585 28373 32597 28376
rect 32631 28373 32643 28407
rect 32585 28367 32643 28373
rect 35526 28364 35532 28416
rect 35584 28404 35590 28416
rect 35897 28407 35955 28413
rect 35897 28404 35909 28407
rect 35584 28376 35909 28404
rect 35584 28364 35590 28376
rect 35897 28373 35909 28376
rect 35943 28373 35955 28407
rect 35897 28367 35955 28373
rect 36262 28364 36268 28416
rect 36320 28404 36326 28416
rect 36357 28407 36415 28413
rect 36357 28404 36369 28407
rect 36320 28376 36369 28404
rect 36320 28364 36326 28376
rect 36357 28373 36369 28376
rect 36403 28373 36415 28407
rect 42334 28404 42340 28416
rect 42295 28376 42340 28404
rect 36357 28367 36415 28373
rect 42334 28364 42340 28376
rect 42392 28364 42398 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 12986 28160 12992 28212
rect 13044 28200 13050 28212
rect 13044 28172 32720 28200
rect 13044 28160 13050 28172
rect 23382 28092 23388 28144
rect 23440 28132 23446 28144
rect 24857 28135 24915 28141
rect 24857 28132 24869 28135
rect 23440 28104 24869 28132
rect 23440 28092 23446 28104
rect 24857 28101 24869 28104
rect 24903 28101 24915 28135
rect 24857 28095 24915 28101
rect 24946 28092 24952 28144
rect 25004 28132 25010 28144
rect 25073 28135 25131 28141
rect 25073 28132 25085 28135
rect 25004 28104 25085 28132
rect 25004 28092 25010 28104
rect 25073 28101 25085 28104
rect 25119 28132 25131 28135
rect 25590 28132 25596 28144
rect 25119 28104 25596 28132
rect 25119 28101 25131 28104
rect 25073 28095 25131 28101
rect 25590 28092 25596 28104
rect 25648 28092 25654 28144
rect 26237 28135 26295 28141
rect 26237 28101 26249 28135
rect 26283 28132 26295 28135
rect 26326 28132 26332 28144
rect 26283 28104 26332 28132
rect 26283 28101 26295 28104
rect 26237 28095 26295 28101
rect 26326 28092 26332 28104
rect 26384 28092 26390 28144
rect 26602 28132 26608 28144
rect 26563 28104 26608 28132
rect 26602 28092 26608 28104
rect 26660 28092 26666 28144
rect 32585 28135 32643 28141
rect 32585 28101 32597 28135
rect 32631 28101 32643 28135
rect 32692 28132 32720 28172
rect 32950 28160 32956 28212
rect 33008 28200 33014 28212
rect 33137 28203 33195 28209
rect 33137 28200 33149 28203
rect 33008 28172 33149 28200
rect 33008 28160 33014 28172
rect 33137 28169 33149 28172
rect 33183 28169 33195 28203
rect 38010 28200 38016 28212
rect 37971 28172 38016 28200
rect 33137 28163 33195 28169
rect 38010 28160 38016 28172
rect 38068 28160 38074 28212
rect 38930 28200 38936 28212
rect 38120 28172 38936 28200
rect 36354 28132 36360 28144
rect 32692 28104 35204 28132
rect 32585 28095 32643 28101
rect 22922 28064 22928 28076
rect 22883 28036 22928 28064
rect 22922 28024 22928 28036
rect 22980 28024 22986 28076
rect 23198 28064 23204 28076
rect 23159 28036 23204 28064
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 23658 28064 23664 28076
rect 23619 28036 23664 28064
rect 23658 28024 23664 28036
rect 23716 28024 23722 28076
rect 23842 28064 23848 28076
rect 23803 28036 23848 28064
rect 23842 28024 23848 28036
rect 23900 28024 23906 28076
rect 24029 28067 24087 28073
rect 24029 28033 24041 28067
rect 24075 28064 24087 28067
rect 24118 28064 24124 28076
rect 24075 28036 24124 28064
rect 24075 28033 24087 28036
rect 24029 28027 24087 28033
rect 24118 28024 24124 28036
rect 24176 28024 24182 28076
rect 24224 28067 24282 28073
rect 24224 28033 24236 28067
rect 24270 28064 24282 28067
rect 24270 28036 24440 28064
rect 24270 28033 24282 28036
rect 24224 28027 24282 28033
rect 23014 27956 23020 28008
rect 23072 27996 23078 28008
rect 23946 27999 24004 28005
rect 23946 27996 23958 27999
rect 23072 27968 23958 27996
rect 23072 27956 23078 27968
rect 23946 27965 23958 27968
rect 23992 27965 24004 27999
rect 23946 27959 24004 27965
rect 22741 27931 22799 27937
rect 22741 27897 22753 27931
rect 22787 27928 22799 27931
rect 23750 27928 23756 27940
rect 22787 27900 23756 27928
rect 22787 27897 22799 27900
rect 22741 27891 22799 27897
rect 23750 27888 23756 27900
rect 23808 27888 23814 27940
rect 24412 27928 24440 28036
rect 26510 28024 26516 28076
rect 26568 28064 26574 28076
rect 28629 28067 28687 28073
rect 28629 28064 28641 28067
rect 26568 28036 28641 28064
rect 26568 28024 26574 28036
rect 28629 28033 28641 28036
rect 28675 28064 28687 28067
rect 29914 28064 29920 28076
rect 28675 28036 29920 28064
rect 28675 28033 28687 28036
rect 28629 28027 28687 28033
rect 29914 28024 29920 28036
rect 29972 28024 29978 28076
rect 30650 28024 30656 28076
rect 30708 28064 30714 28076
rect 30929 28067 30987 28073
rect 30929 28064 30941 28067
rect 30708 28036 30941 28064
rect 30708 28024 30714 28036
rect 30929 28033 30941 28036
rect 30975 28033 30987 28067
rect 32306 28064 32312 28076
rect 32267 28036 32312 28064
rect 30929 28027 30987 28033
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 32600 28064 32628 28095
rect 33045 28067 33103 28073
rect 33045 28064 33057 28067
rect 32600 28036 33057 28064
rect 33045 28033 33057 28036
rect 33091 28033 33103 28067
rect 33045 28027 33103 28033
rect 33229 28067 33287 28073
rect 33229 28033 33241 28067
rect 33275 28033 33287 28067
rect 33229 28027 33287 28033
rect 24486 27956 24492 28008
rect 24544 27996 24550 28008
rect 31205 27999 31263 28005
rect 24544 27968 25360 27996
rect 24544 27956 24550 27968
rect 24762 27928 24768 27940
rect 24412 27900 24768 27928
rect 24762 27888 24768 27900
rect 24820 27888 24826 27940
rect 25222 27928 25228 27940
rect 25183 27900 25228 27928
rect 25222 27888 25228 27900
rect 25280 27888 25286 27940
rect 23109 27863 23167 27869
rect 23109 27829 23121 27863
rect 23155 27860 23167 27863
rect 23474 27860 23480 27872
rect 23155 27832 23480 27860
rect 23155 27829 23167 27832
rect 23109 27823 23167 27829
rect 23474 27820 23480 27832
rect 23532 27820 23538 27872
rect 24397 27863 24455 27869
rect 24397 27829 24409 27863
rect 24443 27860 24455 27863
rect 24854 27860 24860 27872
rect 24443 27832 24860 27860
rect 24443 27829 24455 27832
rect 24397 27823 24455 27829
rect 24854 27820 24860 27832
rect 24912 27820 24918 27872
rect 25041 27863 25099 27869
rect 25041 27829 25053 27863
rect 25087 27860 25099 27863
rect 25332 27860 25360 27968
rect 31205 27965 31217 27999
rect 31251 27996 31263 27999
rect 32582 27996 32588 28008
rect 31251 27968 32588 27996
rect 31251 27965 31263 27968
rect 31205 27959 31263 27965
rect 32582 27956 32588 27968
rect 32640 27956 32646 28008
rect 32674 27956 32680 28008
rect 32732 27996 32738 28008
rect 33244 27996 33272 28027
rect 32732 27968 33272 27996
rect 32732 27956 32738 27968
rect 31021 27931 31079 27937
rect 31021 27897 31033 27931
rect 31067 27928 31079 27931
rect 32692 27928 32720 27956
rect 31067 27900 32720 27928
rect 31067 27897 31079 27900
rect 31021 27891 31079 27897
rect 25087 27832 25360 27860
rect 25087 27829 25099 27832
rect 25041 27823 25099 27829
rect 28534 27820 28540 27872
rect 28592 27860 28598 27872
rect 28721 27863 28779 27869
rect 28721 27860 28733 27863
rect 28592 27832 28733 27860
rect 28592 27820 28598 27832
rect 28721 27829 28733 27832
rect 28767 27829 28779 27863
rect 28721 27823 28779 27829
rect 30374 27820 30380 27872
rect 30432 27860 30438 27872
rect 31113 27863 31171 27869
rect 31113 27860 31125 27863
rect 30432 27832 31125 27860
rect 30432 27820 30438 27832
rect 31113 27829 31125 27832
rect 31159 27829 31171 27863
rect 31113 27823 31171 27829
rect 31938 27820 31944 27872
rect 31996 27860 32002 27872
rect 32401 27863 32459 27869
rect 32401 27860 32413 27863
rect 31996 27832 32413 27860
rect 31996 27820 32002 27832
rect 32401 27829 32413 27832
rect 32447 27829 32459 27863
rect 32401 27823 32459 27829
rect 34790 27820 34796 27872
rect 34848 27860 34854 27872
rect 35069 27863 35127 27869
rect 35069 27860 35081 27863
rect 34848 27832 35081 27860
rect 34848 27820 34854 27832
rect 35069 27829 35081 27832
rect 35115 27829 35127 27863
rect 35176 27860 35204 28104
rect 35268 28104 36360 28132
rect 35268 28073 35296 28104
rect 36354 28092 36360 28104
rect 36412 28092 36418 28144
rect 38120 28132 38148 28172
rect 38930 28160 38936 28172
rect 38988 28160 38994 28212
rect 39945 28203 40003 28209
rect 39945 28169 39957 28203
rect 39991 28200 40003 28203
rect 40126 28200 40132 28212
rect 39991 28172 40132 28200
rect 39991 28169 40003 28172
rect 39945 28163 40003 28169
rect 40126 28160 40132 28172
rect 40184 28160 40190 28212
rect 41506 28160 41512 28212
rect 41564 28200 41570 28212
rect 42061 28203 42119 28209
rect 42061 28200 42073 28203
rect 41564 28172 42073 28200
rect 41564 28160 41570 28172
rect 42061 28169 42073 28172
rect 42107 28169 42119 28203
rect 42061 28163 42119 28169
rect 45738 28160 45744 28212
rect 45796 28209 45802 28212
rect 45796 28200 45805 28209
rect 47854 28200 47860 28212
rect 45796 28172 45841 28200
rect 47815 28172 47860 28200
rect 45796 28163 45805 28172
rect 45796 28160 45802 28163
rect 47854 28160 47860 28172
rect 47912 28160 47918 28212
rect 37936 28104 38148 28132
rect 35253 28067 35311 28073
rect 35253 28033 35265 28067
rect 35299 28033 35311 28067
rect 35253 28027 35311 28033
rect 35345 28067 35403 28073
rect 35345 28033 35357 28067
rect 35391 28033 35403 28067
rect 35345 28027 35403 28033
rect 35621 28067 35679 28073
rect 35621 28033 35633 28067
rect 35667 28064 35679 28067
rect 35986 28064 35992 28076
rect 35667 28036 35992 28064
rect 35667 28033 35679 28036
rect 35621 28027 35679 28033
rect 35360 27928 35388 28027
rect 35986 28024 35992 28036
rect 36044 28024 36050 28076
rect 37936 28073 37964 28104
rect 38470 28092 38476 28144
rect 38528 28132 38534 28144
rect 40948 28135 41006 28141
rect 38528 28104 40724 28132
rect 38528 28092 38534 28104
rect 37921 28067 37979 28073
rect 37921 28033 37933 28067
rect 37967 28033 37979 28067
rect 37921 28027 37979 28033
rect 38010 28024 38016 28076
rect 38068 28064 38074 28076
rect 38105 28067 38163 28073
rect 38105 28064 38117 28067
rect 38068 28036 38117 28064
rect 38068 28024 38074 28036
rect 38105 28033 38117 28036
rect 38151 28033 38163 28067
rect 38105 28027 38163 28033
rect 38832 28067 38890 28073
rect 38832 28033 38844 28067
rect 38878 28064 38890 28067
rect 39114 28064 39120 28076
rect 38878 28036 39120 28064
rect 38878 28033 38890 28036
rect 38832 28027 38890 28033
rect 39114 28024 39120 28036
rect 39172 28024 39178 28076
rect 40696 28073 40724 28104
rect 40948 28101 40960 28135
rect 40994 28132 41006 28135
rect 42334 28132 42340 28144
rect 40994 28104 42340 28132
rect 40994 28101 41006 28104
rect 40948 28095 41006 28101
rect 42334 28092 42340 28104
rect 42392 28092 42398 28144
rect 45830 28132 45836 28144
rect 42720 28104 43944 28132
rect 45791 28104 45836 28132
rect 40681 28067 40739 28073
rect 40681 28033 40693 28067
rect 40727 28033 40739 28067
rect 40681 28027 40739 28033
rect 35434 27956 35440 28008
rect 35492 27996 35498 28008
rect 35529 27999 35587 28005
rect 35529 27996 35541 27999
rect 35492 27968 35541 27996
rect 35492 27956 35498 27968
rect 35529 27965 35541 27968
rect 35575 27965 35587 27999
rect 35529 27959 35587 27965
rect 38470 27956 38476 28008
rect 38528 27996 38534 28008
rect 38565 27999 38623 28005
rect 38565 27996 38577 27999
rect 38528 27968 38577 27996
rect 38528 27956 38534 27968
rect 38565 27965 38577 27968
rect 38611 27965 38623 27999
rect 38565 27959 38623 27965
rect 35618 27928 35624 27940
rect 35360 27900 35624 27928
rect 35618 27888 35624 27900
rect 35676 27888 35682 27940
rect 42720 27860 42748 28104
rect 43162 28073 43168 28076
rect 43156 28027 43168 28073
rect 43220 28064 43226 28076
rect 43220 28036 43256 28064
rect 43162 28024 43168 28027
rect 43220 28024 43226 28036
rect 42886 27996 42892 28008
rect 42847 27968 42892 27996
rect 42886 27956 42892 27968
rect 42944 27956 42950 28008
rect 43916 27996 43944 28104
rect 45830 28092 45836 28104
rect 45888 28092 45894 28144
rect 45940 28104 46612 28132
rect 45940 28076 45968 28104
rect 45649 28067 45707 28073
rect 45649 28033 45661 28067
rect 45695 28064 45707 28067
rect 45738 28064 45744 28076
rect 45695 28036 45744 28064
rect 45695 28033 45707 28036
rect 45649 28027 45707 28033
rect 45738 28024 45744 28036
rect 45796 28024 45802 28076
rect 45922 28024 45928 28076
rect 45980 28064 45986 28076
rect 46385 28067 46443 28073
rect 45980 28036 46025 28064
rect 45980 28024 45986 28036
rect 46385 28033 46397 28067
rect 46431 28064 46443 28067
rect 46474 28064 46480 28076
rect 46431 28036 46480 28064
rect 46431 28033 46443 28036
rect 46385 28027 46443 28033
rect 46474 28024 46480 28036
rect 46532 28024 46538 28076
rect 46584 28073 46612 28104
rect 46569 28067 46627 28073
rect 46569 28033 46581 28067
rect 46615 28033 46627 28067
rect 46569 28027 46627 28033
rect 47486 28024 47492 28076
rect 47544 28064 47550 28076
rect 47765 28067 47823 28073
rect 47765 28064 47777 28067
rect 47544 28036 47777 28064
rect 47544 28024 47550 28036
rect 47765 28033 47777 28036
rect 47811 28033 47823 28067
rect 47765 28027 47823 28033
rect 47504 27996 47532 28024
rect 43916 27968 47532 27996
rect 35176 27832 42748 27860
rect 35069 27823 35127 27829
rect 43806 27820 43812 27872
rect 43864 27860 43870 27872
rect 44269 27863 44327 27869
rect 44269 27860 44281 27863
rect 43864 27832 44281 27860
rect 43864 27820 43870 27832
rect 44269 27829 44281 27832
rect 44315 27829 44327 27863
rect 46382 27860 46388 27872
rect 46343 27832 46388 27860
rect 44269 27823 44327 27829
rect 46382 27820 46388 27832
rect 46440 27820 46446 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 22922 27616 22928 27668
rect 22980 27656 22986 27668
rect 26602 27656 26608 27668
rect 22980 27628 26608 27656
rect 22980 27616 22986 27628
rect 26602 27616 26608 27628
rect 26660 27616 26666 27668
rect 39114 27656 39120 27668
rect 39075 27628 39120 27656
rect 39114 27616 39120 27628
rect 39172 27616 39178 27668
rect 40218 27656 40224 27668
rect 40179 27628 40224 27656
rect 40218 27616 40224 27628
rect 40276 27616 40282 27668
rect 40405 27659 40463 27665
rect 40405 27625 40417 27659
rect 40451 27656 40463 27659
rect 41598 27656 41604 27668
rect 40451 27628 41604 27656
rect 40451 27625 40463 27628
rect 40405 27619 40463 27625
rect 22741 27591 22799 27597
rect 22741 27557 22753 27591
rect 22787 27588 22799 27591
rect 23014 27588 23020 27600
rect 22787 27560 23020 27588
rect 22787 27557 22799 27560
rect 22741 27551 22799 27557
rect 23014 27548 23020 27560
rect 23072 27548 23078 27600
rect 24578 27548 24584 27600
rect 24636 27548 24642 27600
rect 25590 27548 25596 27600
rect 25648 27588 25654 27600
rect 26973 27591 27031 27597
rect 26973 27588 26985 27591
rect 25648 27560 26985 27588
rect 25648 27548 25654 27560
rect 26973 27557 26985 27560
rect 27019 27557 27031 27591
rect 26973 27551 27031 27557
rect 32125 27591 32183 27597
rect 32125 27557 32137 27591
rect 32171 27588 32183 27591
rect 32674 27588 32680 27600
rect 32171 27560 32680 27588
rect 32171 27557 32183 27560
rect 32125 27551 32183 27557
rect 32674 27548 32680 27560
rect 32732 27548 32738 27600
rect 33778 27548 33784 27600
rect 33836 27588 33842 27600
rect 38010 27588 38016 27600
rect 33836 27560 38016 27588
rect 33836 27548 33842 27560
rect 38010 27548 38016 27560
rect 38068 27548 38074 27600
rect 39206 27588 39212 27600
rect 39167 27560 39212 27588
rect 39206 27548 39212 27560
rect 39264 27548 39270 27600
rect 40310 27588 40316 27600
rect 40144 27560 40316 27588
rect 23566 27520 23572 27532
rect 23527 27492 23572 27520
rect 23566 27480 23572 27492
rect 23624 27480 23630 27532
rect 23750 27520 23756 27532
rect 23711 27492 23756 27520
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 24596 27520 24624 27548
rect 24320 27492 24624 27520
rect 22646 27452 22652 27464
rect 22607 27424 22652 27452
rect 22646 27412 22652 27424
rect 22704 27412 22710 27464
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 23106 27452 23112 27464
rect 22879 27424 23112 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 23106 27412 23112 27424
rect 23164 27412 23170 27464
rect 23477 27455 23535 27461
rect 23477 27421 23489 27455
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 23661 27455 23719 27461
rect 23661 27421 23673 27455
rect 23707 27452 23719 27455
rect 24320 27452 24348 27492
rect 26326 27480 26332 27532
rect 26384 27520 26390 27532
rect 26513 27523 26571 27529
rect 26513 27520 26525 27523
rect 26384 27492 26525 27520
rect 26384 27480 26390 27492
rect 26513 27489 26525 27492
rect 26559 27489 26571 27523
rect 26513 27483 26571 27489
rect 29822 27480 29828 27532
rect 29880 27520 29886 27532
rect 29917 27523 29975 27529
rect 29917 27520 29929 27523
rect 29880 27492 29929 27520
rect 29880 27480 29886 27492
rect 29917 27489 29929 27492
rect 29963 27489 29975 27523
rect 29917 27483 29975 27489
rect 31757 27523 31815 27529
rect 31757 27489 31769 27523
rect 31803 27520 31815 27523
rect 31846 27520 31852 27532
rect 31803 27492 31852 27520
rect 31803 27489 31815 27492
rect 31757 27483 31815 27489
rect 31846 27480 31852 27492
rect 31904 27520 31910 27532
rect 32306 27520 32312 27532
rect 31904 27492 32312 27520
rect 31904 27480 31910 27492
rect 32306 27480 32312 27492
rect 32364 27480 32370 27532
rect 35526 27520 35532 27532
rect 35084 27492 35532 27520
rect 23707 27424 24348 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 23492 27384 23520 27415
rect 24394 27412 24400 27464
rect 24452 27452 24458 27464
rect 24854 27461 24860 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24452 27424 24593 27452
rect 24452 27412 24458 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24848 27452 24860 27461
rect 24815 27424 24860 27452
rect 24581 27415 24639 27421
rect 24848 27415 24860 27424
rect 24854 27412 24860 27415
rect 24912 27412 24918 27464
rect 26602 27452 26608 27464
rect 26563 27424 26608 27452
rect 26602 27412 26608 27424
rect 26660 27412 26666 27464
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27433 27415 27491 27421
rect 25590 27384 25596 27396
rect 23492 27356 25596 27384
rect 25590 27344 25596 27356
rect 25648 27344 25654 27396
rect 25682 27344 25688 27396
rect 25740 27384 25746 27396
rect 27448 27384 27476 27415
rect 27522 27412 27528 27464
rect 27580 27452 27586 27464
rect 28077 27455 28135 27461
rect 28077 27452 28089 27455
rect 27580 27424 28089 27452
rect 27580 27412 27586 27424
rect 28077 27421 28089 27424
rect 28123 27421 28135 27455
rect 31938 27452 31944 27464
rect 31899 27424 31944 27452
rect 28077 27415 28135 27421
rect 31938 27412 31944 27424
rect 31996 27412 32002 27464
rect 35084 27461 35112 27492
rect 35526 27480 35532 27492
rect 35584 27480 35590 27532
rect 38028 27520 38056 27548
rect 39393 27523 39451 27529
rect 40144 27528 40172 27560
rect 40310 27548 40316 27560
rect 40368 27548 40374 27600
rect 39393 27520 39405 27523
rect 38028 27492 39405 27520
rect 39393 27489 39405 27492
rect 39439 27520 39451 27523
rect 40052 27520 40172 27528
rect 40420 27520 40448 27619
rect 41598 27616 41604 27628
rect 41656 27616 41662 27668
rect 42061 27659 42119 27665
rect 42061 27625 42073 27659
rect 42107 27656 42119 27659
rect 42426 27656 42432 27668
rect 42107 27628 42432 27656
rect 42107 27625 42119 27628
rect 42061 27619 42119 27625
rect 42426 27616 42432 27628
rect 42484 27616 42490 27668
rect 43162 27656 43168 27668
rect 43123 27628 43168 27656
rect 43162 27616 43168 27628
rect 43220 27616 43226 27668
rect 43898 27656 43904 27668
rect 43859 27628 43904 27656
rect 43898 27616 43904 27628
rect 43956 27616 43962 27668
rect 45922 27616 45928 27668
rect 45980 27656 45986 27668
rect 46109 27659 46167 27665
rect 46109 27656 46121 27659
rect 45980 27628 46121 27656
rect 45980 27616 45986 27628
rect 46109 27625 46121 27628
rect 46155 27625 46167 27659
rect 46109 27619 46167 27625
rect 46474 27616 46480 27668
rect 46532 27656 46538 27668
rect 46753 27659 46811 27665
rect 46753 27656 46765 27659
rect 46532 27628 46765 27656
rect 46532 27616 46538 27628
rect 46753 27625 46765 27628
rect 46799 27625 46811 27659
rect 46753 27619 46811 27625
rect 42886 27548 42892 27600
rect 42944 27588 42950 27600
rect 43254 27588 43260 27600
rect 42944 27560 43260 27588
rect 42944 27548 42950 27560
rect 43254 27548 43260 27560
rect 43312 27588 43318 27600
rect 45554 27588 45560 27600
rect 43312 27560 45560 27588
rect 43312 27548 43318 27560
rect 45554 27548 45560 27560
rect 45612 27548 45618 27600
rect 45756 27560 46796 27588
rect 39439 27500 40172 27520
rect 39439 27492 40080 27500
rect 40236 27492 40448 27520
rect 39439 27489 39451 27492
rect 39393 27483 39451 27489
rect 35069 27455 35127 27461
rect 35069 27421 35081 27455
rect 35115 27421 35127 27455
rect 35342 27452 35348 27464
rect 35303 27424 35348 27452
rect 35069 27415 35127 27421
rect 35342 27412 35348 27424
rect 35400 27412 35406 27464
rect 40236 27462 40264 27492
rect 41506 27480 41512 27532
rect 41564 27520 41570 27532
rect 41693 27523 41751 27529
rect 41693 27520 41705 27523
rect 41564 27492 41705 27520
rect 41564 27480 41570 27492
rect 41693 27489 41705 27492
rect 41739 27489 41751 27523
rect 41693 27483 41751 27489
rect 42996 27492 44128 27520
rect 39117 27455 39175 27461
rect 39117 27421 39129 27455
rect 39163 27452 39175 27455
rect 40160 27452 40264 27462
rect 39163 27434 40264 27452
rect 39163 27424 40188 27434
rect 39163 27421 39175 27424
rect 39117 27415 39175 27421
rect 40310 27412 40316 27464
rect 40368 27412 40374 27464
rect 41598 27412 41604 27464
rect 41656 27452 41662 27464
rect 42996 27461 43024 27492
rect 41877 27455 41935 27461
rect 41877 27452 41889 27455
rect 41656 27424 41889 27452
rect 41656 27412 41662 27424
rect 41877 27421 41889 27424
rect 41923 27421 41935 27455
rect 41877 27415 41935 27421
rect 42981 27455 43039 27461
rect 42981 27421 42993 27455
rect 43027 27421 43039 27455
rect 42981 27415 43039 27421
rect 43073 27455 43131 27461
rect 43073 27421 43085 27455
rect 43119 27452 43131 27455
rect 43346 27452 43352 27464
rect 43119 27424 43352 27452
rect 43119 27421 43131 27424
rect 43073 27415 43131 27421
rect 43346 27412 43352 27424
rect 43404 27412 43410 27464
rect 30190 27393 30196 27396
rect 25740 27356 27476 27384
rect 25740 27344 25746 27356
rect 30184 27347 30196 27393
rect 30248 27384 30254 27396
rect 33686 27384 33692 27396
rect 30248 27356 30284 27384
rect 33647 27356 33692 27384
rect 30190 27344 30196 27347
rect 30248 27344 30254 27356
rect 33686 27344 33692 27356
rect 33744 27344 33750 27396
rect 34885 27387 34943 27393
rect 34885 27353 34897 27387
rect 34931 27384 34943 27387
rect 35894 27384 35900 27396
rect 34931 27356 35900 27384
rect 34931 27353 34943 27356
rect 34885 27347 34943 27353
rect 35894 27344 35900 27356
rect 35952 27344 35958 27396
rect 40037 27387 40095 27393
rect 40037 27353 40049 27387
rect 40083 27384 40095 27387
rect 40126 27384 40132 27396
rect 40083 27356 40132 27384
rect 40083 27353 40095 27356
rect 40037 27347 40095 27353
rect 40126 27344 40132 27356
rect 40184 27344 40190 27396
rect 40328 27384 40356 27412
rect 41046 27384 41052 27396
rect 40328 27356 41052 27384
rect 41046 27344 41052 27356
rect 41104 27384 41110 27396
rect 43257 27387 43315 27393
rect 43257 27384 43269 27387
rect 41104 27356 43269 27384
rect 41104 27344 41110 27356
rect 43257 27353 43269 27356
rect 43303 27353 43315 27387
rect 43714 27384 43720 27396
rect 43675 27356 43720 27384
rect 43257 27347 43315 27353
rect 43714 27344 43720 27356
rect 43772 27344 43778 27396
rect 23290 27316 23296 27328
rect 23251 27288 23296 27316
rect 23290 27276 23296 27288
rect 23348 27276 23354 27328
rect 25958 27316 25964 27328
rect 25919 27288 25964 27316
rect 25958 27276 25964 27288
rect 26016 27276 26022 27328
rect 27525 27319 27583 27325
rect 27525 27285 27537 27319
rect 27571 27316 27583 27319
rect 27614 27316 27620 27328
rect 27571 27288 27620 27316
rect 27571 27285 27583 27288
rect 27525 27279 27583 27285
rect 27614 27276 27620 27288
rect 27672 27276 27678 27328
rect 28166 27316 28172 27328
rect 28127 27288 28172 27316
rect 28166 27276 28172 27288
rect 28224 27276 28230 27328
rect 30650 27276 30656 27328
rect 30708 27316 30714 27328
rect 31297 27319 31355 27325
rect 31297 27316 31309 27319
rect 30708 27288 31309 27316
rect 30708 27276 30714 27288
rect 31297 27285 31309 27288
rect 31343 27285 31355 27319
rect 33778 27316 33784 27328
rect 33739 27288 33784 27316
rect 31297 27279 31355 27285
rect 33778 27276 33784 27288
rect 33836 27276 33842 27328
rect 35253 27319 35311 27325
rect 35253 27285 35265 27319
rect 35299 27316 35311 27319
rect 35342 27316 35348 27328
rect 35299 27288 35348 27316
rect 35299 27285 35311 27288
rect 35253 27279 35311 27285
rect 35342 27276 35348 27288
rect 35400 27276 35406 27328
rect 40237 27319 40295 27325
rect 40237 27285 40249 27319
rect 40283 27316 40295 27319
rect 40402 27316 40408 27328
rect 40283 27288 40408 27316
rect 40283 27285 40295 27288
rect 40237 27279 40295 27285
rect 40402 27276 40408 27288
rect 40460 27276 40466 27328
rect 42426 27276 42432 27328
rect 42484 27316 42490 27328
rect 43622 27316 43628 27328
rect 42484 27288 43628 27316
rect 42484 27276 42490 27288
rect 43622 27276 43628 27288
rect 43680 27316 43686 27328
rect 44100 27325 44128 27492
rect 45646 27480 45652 27532
rect 45704 27520 45710 27532
rect 45756 27529 45784 27560
rect 45741 27523 45799 27529
rect 45741 27520 45753 27523
rect 45704 27492 45753 27520
rect 45704 27480 45710 27492
rect 45741 27489 45753 27492
rect 45787 27489 45799 27523
rect 46661 27523 46719 27529
rect 46661 27520 46673 27523
rect 45741 27483 45799 27489
rect 45940 27492 46673 27520
rect 45940 27461 45968 27492
rect 46661 27489 46673 27492
rect 46707 27489 46719 27523
rect 46661 27483 46719 27489
rect 46768 27464 46796 27560
rect 46842 27480 46848 27532
rect 46900 27520 46906 27532
rect 46900 27492 46945 27520
rect 46900 27480 46906 27492
rect 45925 27455 45983 27461
rect 45925 27421 45937 27455
rect 45971 27421 45983 27455
rect 45925 27415 45983 27421
rect 46569 27455 46627 27461
rect 46569 27421 46581 27455
rect 46615 27452 46627 27455
rect 46750 27452 46756 27464
rect 46615 27424 46756 27452
rect 46615 27421 46627 27424
rect 46569 27415 46627 27421
rect 43917 27319 43975 27325
rect 43917 27316 43929 27319
rect 43680 27288 43929 27316
rect 43680 27276 43686 27288
rect 43917 27285 43929 27288
rect 43963 27285 43975 27319
rect 43917 27279 43975 27285
rect 44085 27319 44143 27325
rect 44085 27285 44097 27319
rect 44131 27316 44143 27319
rect 45940 27316 45968 27415
rect 46750 27412 46756 27424
rect 46808 27412 46814 27464
rect 44131 27288 45968 27316
rect 44131 27285 44143 27288
rect 44085 27279 44143 27285
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 23382 27112 23388 27124
rect 23343 27084 23388 27112
rect 23382 27072 23388 27084
rect 23440 27072 23446 27124
rect 25317 27115 25375 27121
rect 25317 27081 25329 27115
rect 25363 27112 25375 27115
rect 26602 27112 26608 27124
rect 25363 27084 26608 27112
rect 25363 27081 25375 27084
rect 25317 27075 25375 27081
rect 26602 27072 26608 27084
rect 26660 27112 26666 27124
rect 30101 27115 30159 27121
rect 26660 27084 27568 27112
rect 26660 27072 26666 27084
rect 25682 27044 25688 27056
rect 24136 27016 25688 27044
rect 22922 26936 22928 26988
rect 22980 26976 22986 26988
rect 23293 26979 23351 26985
rect 23293 26976 23305 26979
rect 22980 26948 23305 26976
rect 22980 26936 22986 26948
rect 23293 26945 23305 26948
rect 23339 26945 23351 26979
rect 23293 26939 23351 26945
rect 23474 26936 23480 26988
rect 23532 26976 23538 26988
rect 24136 26976 24164 27016
rect 25682 27004 25688 27016
rect 25740 27004 25746 27056
rect 27540 27044 27568 27084
rect 30101 27081 30113 27115
rect 30147 27112 30159 27115
rect 30190 27112 30196 27124
rect 30147 27084 30196 27112
rect 30147 27081 30159 27084
rect 30101 27075 30159 27081
rect 30190 27072 30196 27084
rect 30248 27072 30254 27124
rect 31018 27112 31024 27124
rect 30484 27084 31024 27112
rect 30374 27044 30380 27056
rect 27540 27016 27844 27044
rect 27816 26988 27844 27016
rect 30024 27016 30380 27044
rect 23532 26948 24164 26976
rect 25225 26979 25283 26985
rect 23532 26936 23538 26948
rect 25225 26945 25237 26979
rect 25271 26976 25283 26979
rect 25958 26976 25964 26988
rect 25271 26948 25964 26976
rect 25271 26945 25283 26948
rect 25225 26939 25283 26945
rect 23198 26868 23204 26920
rect 23256 26908 23262 26920
rect 24762 26908 24768 26920
rect 23256 26880 24768 26908
rect 23256 26868 23262 26880
rect 24762 26868 24768 26880
rect 24820 26908 24826 26920
rect 25240 26908 25268 26939
rect 25958 26936 25964 26948
rect 26016 26936 26022 26988
rect 26053 26979 26111 26985
rect 26053 26945 26065 26979
rect 26099 26976 26111 26979
rect 27430 26976 27436 26988
rect 26099 26948 27292 26976
rect 27391 26948 27436 26976
rect 26099 26945 26111 26948
rect 26053 26939 26111 26945
rect 24820 26880 25268 26908
rect 26145 26911 26203 26917
rect 24820 26868 24826 26880
rect 26145 26877 26157 26911
rect 26191 26908 26203 26911
rect 26326 26908 26332 26920
rect 26191 26880 26332 26908
rect 26191 26877 26203 26880
rect 26145 26871 26203 26877
rect 26326 26868 26332 26880
rect 26384 26868 26390 26920
rect 27264 26908 27292 26948
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 27522 26936 27528 26988
rect 27580 26976 27586 26988
rect 27798 26976 27804 26988
rect 27580 26948 27625 26976
rect 27711 26948 27804 26976
rect 27580 26936 27586 26948
rect 27798 26936 27804 26948
rect 27856 26936 27862 26988
rect 30024 26985 30052 27016
rect 30374 27004 30380 27016
rect 30432 27004 30438 27056
rect 30009 26979 30067 26985
rect 30009 26945 30021 26979
rect 30055 26945 30067 26979
rect 30009 26939 30067 26945
rect 30193 26979 30251 26985
rect 30193 26945 30205 26979
rect 30239 26976 30251 26979
rect 30484 26976 30512 27084
rect 31018 27072 31024 27084
rect 31076 27072 31082 27124
rect 31938 27112 31944 27124
rect 31726 27084 31944 27112
rect 30650 27044 30656 27056
rect 30611 27016 30656 27044
rect 30650 27004 30656 27016
rect 30708 27004 30714 27056
rect 30869 27047 30927 27053
rect 30869 27013 30881 27047
rect 30915 27044 30927 27047
rect 31294 27044 31300 27056
rect 30915 27016 31300 27044
rect 30915 27013 30927 27016
rect 30869 27007 30927 27013
rect 31294 27004 31300 27016
rect 31352 27044 31358 27056
rect 31726 27044 31754 27084
rect 31938 27072 31944 27084
rect 31996 27072 32002 27124
rect 34333 27115 34391 27121
rect 34333 27081 34345 27115
rect 34379 27112 34391 27115
rect 34977 27115 35035 27121
rect 34977 27112 34989 27115
rect 34379 27084 34989 27112
rect 34379 27081 34391 27084
rect 34333 27075 34391 27081
rect 34977 27081 34989 27084
rect 35023 27112 35035 27115
rect 35342 27112 35348 27124
rect 35023 27084 35348 27112
rect 35023 27081 35035 27084
rect 34977 27075 35035 27081
rect 35342 27072 35348 27084
rect 35400 27072 35406 27124
rect 36906 27112 36912 27124
rect 36867 27084 36912 27112
rect 36906 27072 36912 27084
rect 36964 27072 36970 27124
rect 43533 27115 43591 27121
rect 43533 27081 43545 27115
rect 43579 27112 43591 27115
rect 43898 27112 43904 27124
rect 43579 27084 43904 27112
rect 43579 27081 43591 27084
rect 43533 27075 43591 27081
rect 43898 27072 43904 27084
rect 43956 27072 43962 27124
rect 46750 27072 46756 27124
rect 46808 27112 46814 27124
rect 47213 27115 47271 27121
rect 47213 27112 47225 27115
rect 46808 27084 47225 27112
rect 46808 27072 46814 27084
rect 47213 27081 47225 27084
rect 47259 27081 47271 27115
rect 47213 27075 47271 27081
rect 38286 27044 38292 27056
rect 31352 27016 31754 27044
rect 32968 27016 35572 27044
rect 31352 27004 31358 27016
rect 30239 26948 30512 26976
rect 30239 26945 30251 26948
rect 30193 26939 30251 26945
rect 27540 26908 27568 26936
rect 32968 26920 32996 27016
rect 33220 26979 33278 26985
rect 33220 26945 33232 26979
rect 33266 26976 33278 26979
rect 33502 26976 33508 26988
rect 33266 26948 33508 26976
rect 33266 26945 33278 26948
rect 33220 26939 33278 26945
rect 33502 26936 33508 26948
rect 33560 26936 33566 26988
rect 33686 26936 33692 26988
rect 33744 26976 33750 26988
rect 34793 26979 34851 26985
rect 34793 26976 34805 26979
rect 33744 26948 34805 26976
rect 33744 26936 33750 26948
rect 34793 26945 34805 26948
rect 34839 26945 34851 26979
rect 35066 26976 35072 26988
rect 35027 26948 35072 26976
rect 34793 26939 34851 26945
rect 32950 26908 32956 26920
rect 27264 26880 27568 26908
rect 32911 26880 32956 26908
rect 32950 26868 32956 26880
rect 33008 26868 33014 26920
rect 34808 26908 34836 26939
rect 35066 26936 35072 26948
rect 35124 26936 35130 26988
rect 35544 26985 35572 27016
rect 35636 27016 38292 27044
rect 35529 26979 35587 26985
rect 35529 26945 35541 26979
rect 35575 26945 35587 26979
rect 35529 26939 35587 26945
rect 35636 26908 35664 27016
rect 38286 27004 38292 27016
rect 38344 27004 38350 27056
rect 43349 27047 43407 27053
rect 43349 27013 43361 27047
rect 43395 27044 43407 27047
rect 43714 27044 43720 27056
rect 43395 27016 43720 27044
rect 43395 27013 43407 27016
rect 43349 27007 43407 27013
rect 43714 27004 43720 27016
rect 43772 27004 43778 27056
rect 46100 27047 46158 27053
rect 46100 27013 46112 27047
rect 46146 27044 46158 27047
rect 46382 27044 46388 27056
rect 46146 27016 46388 27044
rect 46146 27013 46158 27016
rect 46100 27007 46158 27013
rect 46382 27004 46388 27016
rect 46440 27004 46446 27056
rect 35796 26979 35854 26985
rect 35796 26945 35808 26979
rect 35842 26976 35854 26979
rect 36170 26976 36176 26988
rect 35842 26948 36176 26976
rect 35842 26945 35854 26948
rect 35796 26939 35854 26945
rect 36170 26936 36176 26948
rect 36228 26936 36234 26988
rect 43622 26976 43628 26988
rect 43583 26948 43628 26976
rect 43622 26936 43628 26948
rect 43680 26936 43686 26988
rect 45554 26936 45560 26988
rect 45612 26976 45618 26988
rect 45833 26979 45891 26985
rect 45833 26976 45845 26979
rect 45612 26948 45845 26976
rect 45612 26936 45618 26948
rect 45833 26945 45845 26948
rect 45879 26945 45891 26979
rect 45833 26939 45891 26945
rect 46934 26936 46940 26988
rect 46992 26976 46998 26988
rect 47578 26976 47584 26988
rect 46992 26948 47584 26976
rect 46992 26936 46998 26948
rect 47578 26936 47584 26948
rect 47636 26976 47642 26988
rect 47765 26979 47823 26985
rect 47765 26976 47777 26979
rect 47636 26948 47777 26976
rect 47636 26936 47642 26948
rect 47765 26945 47777 26948
rect 47811 26945 47823 26979
rect 47765 26939 47823 26945
rect 34808 26880 35664 26908
rect 27338 26800 27344 26852
rect 27396 26840 27402 26852
rect 30650 26840 30656 26852
rect 27396 26812 30656 26840
rect 27396 26800 27402 26812
rect 30650 26800 30656 26812
rect 30708 26800 30714 26852
rect 31846 26840 31852 26852
rect 30852 26812 31852 26840
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 24670 26772 24676 26784
rect 23624 26744 24676 26772
rect 23624 26732 23630 26744
rect 24670 26732 24676 26744
rect 24728 26772 24734 26784
rect 26329 26775 26387 26781
rect 26329 26772 26341 26775
rect 24728 26744 26341 26772
rect 24728 26732 24734 26744
rect 26329 26741 26341 26744
rect 26375 26741 26387 26775
rect 26329 26735 26387 26741
rect 27249 26775 27307 26781
rect 27249 26741 27261 26775
rect 27295 26772 27307 26775
rect 27430 26772 27436 26784
rect 27295 26744 27436 26772
rect 27295 26741 27307 26744
rect 27249 26735 27307 26741
rect 27430 26732 27436 26744
rect 27488 26732 27494 26784
rect 27706 26772 27712 26784
rect 27619 26744 27712 26772
rect 27706 26732 27712 26744
rect 27764 26772 27770 26784
rect 30852 26781 30880 26812
rect 31846 26800 31852 26812
rect 31904 26800 31910 26852
rect 36722 26800 36728 26852
rect 36780 26840 36786 26852
rect 37182 26840 37188 26852
rect 36780 26812 37188 26840
rect 36780 26800 36786 26812
rect 37182 26800 37188 26812
rect 37240 26840 37246 26852
rect 41598 26840 41604 26852
rect 37240 26812 41604 26840
rect 37240 26800 37246 26812
rect 41598 26800 41604 26812
rect 41656 26800 41662 26852
rect 43346 26840 43352 26852
rect 43307 26812 43352 26840
rect 43346 26800 43352 26812
rect 43404 26800 43410 26852
rect 30837 26775 30895 26781
rect 30837 26772 30849 26775
rect 27764 26744 30849 26772
rect 27764 26732 27770 26744
rect 30837 26741 30849 26744
rect 30883 26741 30895 26775
rect 34790 26772 34796 26784
rect 34751 26744 34796 26772
rect 30837 26735 30895 26741
rect 34790 26732 34796 26744
rect 34848 26732 34854 26784
rect 35066 26732 35072 26784
rect 35124 26772 35130 26784
rect 37826 26772 37832 26784
rect 35124 26744 37832 26772
rect 35124 26732 35130 26744
rect 37826 26732 37832 26744
rect 37884 26732 37890 26784
rect 38286 26732 38292 26784
rect 38344 26772 38350 26784
rect 45646 26772 45652 26784
rect 38344 26744 45652 26772
rect 38344 26732 38350 26744
rect 45646 26732 45652 26744
rect 45704 26732 45710 26784
rect 47854 26772 47860 26784
rect 47815 26744 47860 26772
rect 47854 26732 47860 26744
rect 47912 26732 47918 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 31754 26528 31760 26580
rect 31812 26568 31818 26580
rect 32493 26571 32551 26577
rect 32493 26568 32505 26571
rect 31812 26540 32505 26568
rect 31812 26528 31818 26540
rect 32493 26537 32505 26540
rect 32539 26568 32551 26571
rect 32950 26568 32956 26580
rect 32539 26540 32956 26568
rect 32539 26537 32551 26540
rect 32493 26531 32551 26537
rect 32950 26528 32956 26540
rect 33008 26528 33014 26580
rect 33502 26568 33508 26580
rect 33463 26540 33508 26568
rect 33502 26528 33508 26540
rect 33560 26528 33566 26580
rect 33873 26571 33931 26577
rect 33873 26537 33885 26571
rect 33919 26568 33931 26571
rect 36538 26568 36544 26580
rect 33919 26540 36544 26568
rect 33919 26537 33931 26540
rect 33873 26531 33931 26537
rect 36538 26528 36544 26540
rect 36596 26528 36602 26580
rect 39482 26528 39488 26580
rect 39540 26568 39546 26580
rect 40402 26568 40408 26580
rect 39540 26540 40408 26568
rect 39540 26528 39546 26540
rect 40402 26528 40408 26540
rect 40460 26528 40466 26580
rect 43622 26528 43628 26580
rect 43680 26568 43686 26580
rect 43809 26571 43867 26577
rect 43809 26568 43821 26571
rect 43680 26540 43821 26568
rect 43680 26528 43686 26540
rect 43809 26537 43821 26540
rect 43855 26568 43867 26571
rect 43855 26540 44588 26568
rect 43855 26537 43867 26540
rect 43809 26531 43867 26537
rect 35713 26503 35771 26509
rect 35713 26469 35725 26503
rect 35759 26500 35771 26503
rect 37182 26500 37188 26512
rect 35759 26472 37188 26500
rect 35759 26469 35771 26472
rect 35713 26463 35771 26469
rect 37182 26460 37188 26472
rect 37240 26460 37246 26512
rect 39209 26503 39267 26509
rect 39209 26469 39221 26503
rect 39255 26469 39267 26503
rect 39209 26463 39267 26469
rect 28074 26432 28080 26444
rect 27356 26404 28080 26432
rect 26326 26364 26332 26376
rect 26287 26336 26332 26364
rect 26326 26324 26332 26336
rect 26384 26324 26390 26376
rect 27356 26373 27384 26404
rect 28074 26392 28080 26404
rect 28132 26392 28138 26444
rect 34790 26432 34796 26444
rect 33704 26404 34796 26432
rect 26513 26367 26571 26373
rect 26513 26333 26525 26367
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26364 26755 26367
rect 27157 26367 27215 26373
rect 27157 26364 27169 26367
rect 26743 26336 27169 26364
rect 26743 26333 26755 26336
rect 26697 26327 26755 26333
rect 27157 26333 27169 26336
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 27305 26367 27384 26373
rect 27305 26333 27317 26367
rect 27351 26336 27384 26367
rect 27351 26333 27363 26336
rect 27305 26327 27363 26333
rect 26528 26228 26556 26327
rect 27430 26324 27436 26376
rect 27488 26364 27494 26376
rect 27706 26373 27712 26376
rect 27663 26367 27712 26373
rect 27488 26336 27533 26364
rect 27488 26324 27494 26336
rect 27663 26333 27675 26367
rect 27709 26333 27712 26367
rect 27663 26327 27712 26333
rect 27706 26324 27712 26327
rect 27764 26324 27770 26376
rect 27798 26324 27804 26376
rect 27856 26324 27862 26376
rect 33704 26373 33732 26404
rect 34790 26392 34796 26404
rect 34848 26392 34854 26444
rect 35434 26432 35440 26444
rect 35395 26404 35440 26432
rect 35434 26392 35440 26404
rect 35492 26392 35498 26444
rect 39224 26432 39252 26463
rect 40218 26460 40224 26512
rect 40276 26500 40282 26512
rect 44361 26503 44419 26509
rect 40276 26472 40540 26500
rect 40276 26460 40282 26472
rect 40512 26441 40540 26472
rect 44361 26469 44373 26503
rect 44407 26469 44419 26503
rect 44361 26463 44419 26469
rect 40497 26435 40555 26441
rect 39224 26404 40264 26432
rect 33689 26367 33747 26373
rect 33689 26333 33701 26367
rect 33735 26333 33747 26367
rect 33689 26327 33747 26333
rect 33965 26367 34023 26373
rect 33965 26333 33977 26367
rect 34011 26364 34023 26367
rect 35342 26364 35348 26376
rect 34011 26336 35348 26364
rect 34011 26333 34023 26336
rect 33965 26327 34023 26333
rect 35342 26324 35348 26336
rect 35400 26324 35406 26376
rect 38010 26364 38016 26376
rect 37971 26336 38016 26364
rect 38010 26324 38016 26336
rect 38068 26364 38074 26376
rect 38470 26364 38476 26376
rect 38068 26336 38476 26364
rect 38068 26324 38074 26336
rect 38470 26324 38476 26336
rect 38528 26324 38534 26376
rect 39482 26364 39488 26376
rect 39443 26336 39488 26364
rect 39482 26324 39488 26336
rect 39540 26324 39546 26376
rect 40236 26373 40264 26404
rect 40497 26401 40509 26435
rect 40543 26401 40555 26435
rect 44376 26432 44404 26463
rect 40497 26395 40555 26401
rect 43640 26404 44404 26432
rect 44560 26432 44588 26540
rect 46661 26435 46719 26441
rect 44560 26404 44680 26432
rect 43640 26373 43668 26404
rect 40221 26367 40279 26373
rect 40221 26333 40233 26367
rect 40267 26333 40279 26367
rect 40221 26327 40279 26333
rect 43625 26367 43683 26373
rect 43625 26333 43637 26367
rect 43671 26333 43683 26367
rect 43625 26327 43683 26333
rect 43898 26324 43904 26376
rect 43956 26364 43962 26376
rect 44542 26364 44548 26376
rect 43956 26336 44548 26364
rect 43956 26324 43962 26336
rect 44542 26324 44548 26336
rect 44600 26324 44606 26376
rect 44652 26373 44680 26404
rect 46661 26401 46673 26435
rect 46707 26432 46719 26435
rect 47854 26432 47860 26444
rect 46707 26404 47860 26432
rect 46707 26401 46719 26404
rect 46661 26395 46719 26401
rect 47854 26392 47860 26404
rect 47912 26392 47918 26444
rect 48222 26432 48228 26444
rect 48183 26404 48228 26432
rect 48222 26392 48228 26404
rect 48280 26392 48286 26444
rect 44637 26367 44695 26373
rect 44637 26333 44649 26367
rect 44683 26333 44695 26367
rect 44637 26327 44695 26333
rect 46477 26367 46535 26373
rect 46477 26333 46489 26367
rect 46523 26333 46535 26367
rect 46477 26327 46535 26333
rect 27525 26299 27583 26305
rect 27525 26265 27537 26299
rect 27571 26296 27583 26299
rect 27816 26296 27844 26324
rect 31202 26296 31208 26308
rect 27571 26268 27844 26296
rect 31163 26268 31208 26296
rect 27571 26265 27583 26268
rect 27525 26259 27583 26265
rect 31202 26256 31208 26268
rect 31260 26296 31266 26308
rect 36449 26299 36507 26305
rect 36449 26296 36461 26299
rect 31260 26268 36461 26296
rect 31260 26256 31266 26268
rect 36449 26265 36461 26268
rect 36495 26296 36507 26299
rect 36722 26296 36728 26308
rect 36495 26268 36728 26296
rect 36495 26265 36507 26268
rect 36449 26259 36507 26265
rect 36722 26256 36728 26268
rect 36780 26256 36786 26308
rect 36814 26256 36820 26308
rect 36872 26296 36878 26308
rect 36872 26268 38654 26296
rect 36872 26256 36878 26268
rect 38626 26240 38654 26268
rect 38746 26256 38752 26308
rect 38804 26296 38810 26308
rect 39209 26299 39267 26305
rect 39209 26296 39221 26299
rect 38804 26268 39221 26296
rect 38804 26256 38810 26268
rect 39209 26265 39221 26268
rect 39255 26265 39267 26299
rect 39209 26259 39267 26265
rect 39393 26299 39451 26305
rect 39393 26265 39405 26299
rect 39439 26296 39451 26299
rect 44361 26299 44419 26305
rect 39439 26268 40264 26296
rect 39439 26265 39451 26268
rect 39393 26259 39451 26265
rect 40236 26240 40264 26268
rect 44361 26265 44373 26299
rect 44407 26296 44419 26299
rect 45646 26296 45652 26308
rect 44407 26268 45652 26296
rect 44407 26265 44419 26268
rect 44361 26259 44419 26265
rect 45646 26256 45652 26268
rect 45704 26256 45710 26308
rect 46492 26296 46520 26327
rect 47946 26296 47952 26308
rect 46492 26268 47952 26296
rect 47946 26256 47952 26268
rect 48004 26256 48010 26308
rect 27338 26228 27344 26240
rect 26528 26200 27344 26228
rect 27338 26188 27344 26200
rect 27396 26188 27402 26240
rect 27798 26228 27804 26240
rect 27759 26200 27804 26228
rect 27798 26188 27804 26200
rect 27856 26188 27862 26240
rect 32582 26188 32588 26240
rect 32640 26228 32646 26240
rect 37918 26228 37924 26240
rect 32640 26200 37924 26228
rect 32640 26188 32646 26200
rect 37918 26188 37924 26200
rect 37976 26188 37982 26240
rect 38626 26200 38660 26240
rect 38654 26188 38660 26200
rect 38712 26188 38718 26240
rect 40037 26231 40095 26237
rect 40037 26197 40049 26231
rect 40083 26228 40095 26231
rect 40126 26228 40132 26240
rect 40083 26200 40132 26228
rect 40083 26197 40095 26200
rect 40037 26191 40095 26197
rect 40126 26188 40132 26200
rect 40184 26188 40190 26240
rect 40218 26188 40224 26240
rect 40276 26188 40282 26240
rect 43441 26231 43499 26237
rect 43441 26197 43453 26231
rect 43487 26228 43499 26231
rect 43530 26228 43536 26240
rect 43487 26200 43536 26228
rect 43487 26197 43499 26200
rect 43441 26191 43499 26197
rect 43530 26188 43536 26200
rect 43588 26188 43594 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 29822 25984 29828 26036
rect 29880 26024 29886 26036
rect 29917 26027 29975 26033
rect 29917 26024 29929 26027
rect 29880 25996 29929 26024
rect 29880 25984 29886 25996
rect 29917 25993 29929 25996
rect 29963 25993 29975 26027
rect 29917 25987 29975 25993
rect 35434 25984 35440 26036
rect 35492 26024 35498 26036
rect 35621 26027 35679 26033
rect 35621 26024 35633 26027
rect 35492 25996 35633 26024
rect 35492 25984 35498 25996
rect 35621 25993 35633 25996
rect 35667 25993 35679 26027
rect 36170 26024 36176 26036
rect 36131 25996 36176 26024
rect 35621 25987 35679 25993
rect 36170 25984 36176 25996
rect 36228 25984 36234 26036
rect 36538 26024 36544 26036
rect 36451 25996 36544 26024
rect 36538 25984 36544 25996
rect 36596 26024 36602 26036
rect 36596 25996 37688 26024
rect 36596 25984 36602 25996
rect 27798 25956 27804 25968
rect 27172 25928 27804 25956
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25857 22339 25891
rect 22281 25851 22339 25857
rect 22189 25823 22247 25829
rect 22189 25789 22201 25823
rect 22235 25789 22247 25823
rect 22296 25820 22324 25851
rect 23382 25848 23388 25900
rect 23440 25888 23446 25900
rect 27172 25897 27200 25928
rect 27798 25916 27804 25928
rect 27856 25916 27862 25968
rect 28629 25959 28687 25965
rect 28629 25925 28641 25959
rect 28675 25956 28687 25959
rect 31202 25956 31208 25968
rect 28675 25928 31208 25956
rect 28675 25925 28687 25928
rect 28629 25919 28687 25925
rect 31202 25916 31208 25928
rect 31260 25916 31266 25968
rect 32401 25959 32459 25965
rect 32401 25956 32413 25959
rect 31726 25928 32413 25956
rect 24285 25891 24343 25897
rect 24285 25888 24297 25891
rect 23440 25860 24297 25888
rect 23440 25848 23446 25860
rect 24285 25857 24297 25860
rect 24331 25857 24343 25891
rect 24285 25851 24343 25857
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27338 25888 27344 25900
rect 27299 25860 27344 25888
rect 27157 25851 27215 25857
rect 27338 25848 27344 25860
rect 27396 25848 27402 25900
rect 27709 25891 27767 25897
rect 27709 25857 27721 25891
rect 27755 25888 27767 25891
rect 27982 25888 27988 25900
rect 27755 25860 27988 25888
rect 27755 25857 27767 25860
rect 27709 25851 27767 25857
rect 27982 25848 27988 25860
rect 28040 25848 28046 25900
rect 30837 25891 30895 25897
rect 30837 25857 30849 25891
rect 30883 25888 30895 25891
rect 30926 25888 30932 25900
rect 30883 25860 30932 25888
rect 30883 25857 30895 25860
rect 30837 25851 30895 25857
rect 30926 25848 30932 25860
rect 30984 25848 30990 25900
rect 31021 25891 31079 25897
rect 31021 25857 31033 25891
rect 31067 25888 31079 25891
rect 31726 25888 31754 25928
rect 32401 25925 32413 25928
rect 32447 25956 32459 25959
rect 33686 25956 33692 25968
rect 32447 25928 33692 25956
rect 32447 25925 32459 25928
rect 32401 25919 32459 25925
rect 33686 25916 33692 25928
rect 33744 25916 33750 25968
rect 35526 25888 35532 25900
rect 31067 25860 31754 25888
rect 35487 25860 35532 25888
rect 31067 25857 31079 25860
rect 31021 25851 31079 25857
rect 23934 25820 23940 25832
rect 22296 25792 23940 25820
rect 22189 25783 22247 25789
rect 22204 25752 22232 25783
rect 23934 25780 23940 25792
rect 23992 25780 23998 25832
rect 24029 25823 24087 25829
rect 24029 25789 24041 25823
rect 24075 25789 24087 25823
rect 24029 25783 24087 25789
rect 22922 25752 22928 25764
rect 22204 25724 22928 25752
rect 22922 25712 22928 25724
rect 22980 25712 22986 25764
rect 1578 25644 1584 25696
rect 1636 25684 1642 25696
rect 2317 25687 2375 25693
rect 2317 25684 2329 25687
rect 1636 25656 2329 25684
rect 1636 25644 1642 25656
rect 2317 25653 2329 25656
rect 2363 25653 2375 25687
rect 2317 25647 2375 25653
rect 22370 25644 22376 25696
rect 22428 25684 22434 25696
rect 22557 25687 22615 25693
rect 22557 25684 22569 25687
rect 22428 25656 22569 25684
rect 22428 25644 22434 25656
rect 22557 25653 22569 25656
rect 22603 25653 22615 25687
rect 24044 25684 24072 25783
rect 26326 25780 26332 25832
rect 26384 25820 26390 25832
rect 27433 25823 27491 25829
rect 27433 25820 27445 25823
rect 26384 25792 27445 25820
rect 26384 25780 26390 25792
rect 27433 25789 27445 25792
rect 27479 25789 27491 25823
rect 27433 25783 27491 25789
rect 27525 25823 27583 25829
rect 27525 25789 27537 25823
rect 27571 25789 27583 25823
rect 27525 25783 27583 25789
rect 24394 25684 24400 25696
rect 24044 25656 24400 25684
rect 22557 25647 22615 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 25406 25684 25412 25696
rect 25367 25656 25412 25684
rect 25406 25644 25412 25656
rect 25464 25644 25470 25696
rect 27430 25644 27436 25696
rect 27488 25684 27494 25696
rect 27540 25684 27568 25783
rect 30742 25780 30748 25832
rect 30800 25820 30806 25832
rect 31036 25820 31064 25851
rect 35526 25848 35532 25860
rect 35584 25848 35590 25900
rect 35713 25891 35771 25897
rect 35713 25857 35725 25891
rect 35759 25888 35771 25891
rect 36354 25888 36360 25900
rect 35759 25860 36360 25888
rect 35759 25857 35771 25860
rect 35713 25851 35771 25857
rect 36354 25848 36360 25860
rect 36412 25848 36418 25900
rect 36556 25897 36584 25984
rect 37553 25959 37611 25965
rect 37553 25956 37565 25959
rect 36648 25928 37565 25956
rect 36648 25897 36676 25928
rect 37553 25925 37565 25928
rect 37599 25925 37611 25959
rect 37553 25919 37611 25925
rect 36449 25891 36507 25897
rect 36449 25857 36461 25891
rect 36495 25857 36507 25891
rect 36449 25851 36507 25857
rect 36541 25891 36599 25897
rect 36541 25857 36553 25891
rect 36587 25857 36599 25891
rect 36541 25851 36599 25857
rect 36633 25891 36691 25897
rect 36633 25857 36645 25891
rect 36679 25857 36691 25891
rect 36633 25851 36691 25857
rect 30800 25792 31064 25820
rect 36464 25820 36492 25851
rect 36722 25848 36728 25900
rect 36780 25888 36786 25900
rect 36817 25891 36875 25897
rect 36817 25888 36829 25891
rect 36780 25860 36829 25888
rect 36780 25848 36786 25860
rect 36817 25857 36829 25860
rect 36863 25857 36875 25891
rect 36817 25851 36875 25857
rect 37182 25848 37188 25900
rect 37240 25888 37246 25900
rect 37660 25897 37688 25996
rect 40218 25984 40224 26036
rect 40276 26024 40282 26036
rect 40497 26027 40555 26033
rect 40497 26024 40509 26027
rect 40276 25996 40509 26024
rect 40276 25984 40282 25996
rect 40497 25993 40509 25996
rect 40543 25993 40555 26027
rect 40497 25987 40555 25993
rect 44542 25984 44548 26036
rect 44600 26024 44606 26036
rect 44637 26027 44695 26033
rect 44637 26024 44649 26027
rect 44600 25996 44649 26024
rect 44600 25984 44606 25996
rect 44637 25993 44649 25996
rect 44683 25993 44695 26027
rect 44637 25987 44695 25993
rect 47210 25956 47216 25968
rect 39132 25928 41414 25956
rect 47171 25928 47216 25956
rect 37461 25891 37519 25897
rect 37461 25888 37473 25891
rect 37240 25860 37473 25888
rect 37240 25848 37246 25860
rect 37461 25857 37473 25860
rect 37507 25857 37519 25891
rect 37461 25851 37519 25857
rect 37645 25891 37703 25897
rect 37645 25857 37657 25891
rect 37691 25857 37703 25891
rect 37645 25851 37703 25857
rect 36906 25820 36912 25832
rect 36464 25792 36912 25820
rect 30800 25780 30806 25792
rect 36906 25780 36912 25792
rect 36964 25780 36970 25832
rect 37660 25820 37688 25851
rect 37826 25848 37832 25900
rect 37884 25888 37890 25900
rect 39132 25897 39160 25928
rect 38289 25891 38347 25897
rect 38289 25888 38301 25891
rect 37884 25860 38301 25888
rect 37884 25848 37890 25860
rect 38289 25857 38301 25860
rect 38335 25857 38347 25891
rect 38289 25851 38347 25857
rect 39117 25891 39175 25897
rect 39117 25857 39129 25891
rect 39163 25857 39175 25891
rect 39117 25851 39175 25857
rect 39384 25891 39442 25897
rect 39384 25857 39396 25891
rect 39430 25888 39442 25891
rect 40126 25888 40132 25900
rect 39430 25860 40132 25888
rect 39430 25857 39442 25860
rect 39384 25851 39442 25857
rect 40126 25848 40132 25860
rect 40184 25848 40190 25900
rect 41386 25888 41414 25928
rect 47210 25916 47216 25928
rect 47268 25916 47274 25968
rect 43254 25888 43260 25900
rect 41386 25860 43260 25888
rect 43254 25848 43260 25860
rect 43312 25848 43318 25900
rect 43530 25897 43536 25900
rect 43524 25888 43536 25897
rect 43491 25860 43536 25888
rect 43524 25851 43536 25860
rect 43530 25848 43536 25851
rect 43588 25848 43594 25900
rect 47946 25888 47952 25900
rect 47907 25860 47952 25888
rect 47946 25848 47952 25860
rect 48004 25848 48010 25900
rect 45373 25823 45431 25829
rect 37660 25792 38240 25820
rect 38212 25696 38240 25792
rect 45373 25789 45385 25823
rect 45419 25789 45431 25823
rect 45373 25783 45431 25789
rect 45557 25823 45615 25829
rect 45557 25789 45569 25823
rect 45603 25820 45615 25823
rect 47118 25820 47124 25832
rect 45603 25792 47124 25820
rect 45603 25789 45615 25792
rect 45557 25783 45615 25789
rect 45388 25752 45416 25783
rect 47118 25780 47124 25792
rect 47176 25780 47182 25832
rect 46842 25752 46848 25764
rect 45388 25724 46848 25752
rect 46842 25712 46848 25724
rect 46900 25712 46906 25764
rect 27488 25656 27568 25684
rect 27488 25644 27494 25656
rect 27706 25644 27712 25696
rect 27764 25684 27770 25696
rect 27893 25687 27951 25693
rect 27893 25684 27905 25687
rect 27764 25656 27905 25684
rect 27764 25644 27770 25656
rect 27893 25653 27905 25656
rect 27939 25653 27951 25687
rect 30834 25684 30840 25696
rect 30795 25656 30840 25684
rect 27893 25647 27951 25653
rect 30834 25644 30840 25656
rect 30892 25644 30898 25696
rect 32490 25684 32496 25696
rect 32451 25656 32496 25684
rect 32490 25644 32496 25656
rect 32548 25644 32554 25696
rect 38194 25644 38200 25696
rect 38252 25684 38258 25696
rect 38381 25687 38439 25693
rect 38381 25684 38393 25687
rect 38252 25656 38393 25684
rect 38252 25644 38258 25656
rect 38381 25653 38393 25656
rect 38427 25653 38439 25687
rect 38381 25647 38439 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 23382 25480 23388 25492
rect 23343 25452 23388 25480
rect 23382 25440 23388 25452
rect 23440 25440 23446 25492
rect 23934 25440 23940 25492
rect 23992 25480 23998 25492
rect 24673 25483 24731 25489
rect 24673 25480 24685 25483
rect 23992 25452 24685 25480
rect 23992 25440 23998 25452
rect 24673 25449 24685 25452
rect 24719 25480 24731 25483
rect 26326 25480 26332 25492
rect 24719 25452 26332 25480
rect 24719 25449 24731 25452
rect 24673 25443 24731 25449
rect 26326 25440 26332 25452
rect 26384 25440 26390 25492
rect 28074 25480 28080 25492
rect 28035 25452 28080 25480
rect 28074 25440 28080 25452
rect 28132 25440 28138 25492
rect 36354 25480 36360 25492
rect 36315 25452 36360 25480
rect 36354 25440 36360 25452
rect 36412 25440 36418 25492
rect 38749 25415 38807 25421
rect 38749 25381 38761 25415
rect 38795 25412 38807 25415
rect 38838 25412 38844 25424
rect 38795 25384 38844 25412
rect 38795 25381 38807 25384
rect 38749 25375 38807 25381
rect 38838 25372 38844 25384
rect 38896 25372 38902 25424
rect 41417 25415 41475 25421
rect 41417 25381 41429 25415
rect 41463 25412 41475 25415
rect 42242 25412 42248 25424
rect 41463 25384 42248 25412
rect 41463 25381 41475 25384
rect 41417 25375 41475 25381
rect 42242 25372 42248 25384
rect 42300 25372 42306 25424
rect 46014 25372 46020 25424
rect 46072 25372 46078 25424
rect 1578 25344 1584 25356
rect 1539 25316 1584 25344
rect 1578 25304 1584 25316
rect 1636 25304 1642 25356
rect 2774 25344 2780 25356
rect 2735 25316 2780 25344
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 28166 25344 28172 25356
rect 23676 25316 24624 25344
rect 22738 25276 22744 25288
rect 22651 25248 22744 25276
rect 22738 25236 22744 25248
rect 22796 25276 22802 25288
rect 23290 25276 23296 25288
rect 22796 25248 23296 25276
rect 22796 25236 22802 25248
rect 23290 25236 23296 25248
rect 23348 25236 23354 25288
rect 23676 25285 23704 25316
rect 23661 25279 23719 25285
rect 23661 25245 23673 25279
rect 23707 25245 23719 25279
rect 23661 25239 23719 25245
rect 23753 25279 23811 25285
rect 23753 25245 23765 25279
rect 23799 25245 23811 25279
rect 23753 25239 23811 25245
rect 1762 25208 1768 25220
rect 1723 25180 1768 25208
rect 1762 25168 1768 25180
rect 1820 25168 1826 25220
rect 22370 25168 22376 25220
rect 22428 25208 22434 25220
rect 22557 25211 22615 25217
rect 22557 25208 22569 25211
rect 22428 25180 22569 25208
rect 22428 25168 22434 25180
rect 22557 25177 22569 25180
rect 22603 25177 22615 25211
rect 23768 25208 23796 25239
rect 23842 25236 23848 25288
rect 23900 25276 23906 25288
rect 23900 25248 23945 25276
rect 23900 25236 23906 25248
rect 24026 25236 24032 25288
rect 24084 25276 24090 25288
rect 24596 25285 24624 25316
rect 27816 25316 28172 25344
rect 24581 25279 24639 25285
rect 24084 25248 24129 25276
rect 24084 25236 24090 25248
rect 24581 25245 24593 25279
rect 24627 25276 24639 25279
rect 24946 25276 24952 25288
rect 24627 25248 24952 25276
rect 24627 25245 24639 25248
rect 24581 25239 24639 25245
rect 24946 25236 24952 25248
rect 25004 25276 25010 25288
rect 25406 25276 25412 25288
rect 25004 25248 25412 25276
rect 25004 25236 25010 25248
rect 25406 25236 25412 25248
rect 25464 25236 25470 25288
rect 27433 25279 27491 25285
rect 27433 25245 27445 25279
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 27571 25279 27629 25285
rect 27571 25245 27583 25279
rect 27617 25276 27629 25279
rect 27816 25276 27844 25316
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 30926 25304 30932 25356
rect 30984 25344 30990 25356
rect 31665 25347 31723 25353
rect 31665 25344 31677 25347
rect 30984 25316 31677 25344
rect 30984 25304 30990 25316
rect 31665 25313 31677 25316
rect 31711 25313 31723 25347
rect 31665 25307 31723 25313
rect 31849 25347 31907 25353
rect 31849 25313 31861 25347
rect 31895 25344 31907 25347
rect 32582 25344 32588 25356
rect 31895 25316 32588 25344
rect 31895 25313 31907 25316
rect 31849 25307 31907 25313
rect 32582 25304 32588 25316
rect 32640 25304 32646 25356
rect 35342 25304 35348 25356
rect 35400 25344 35406 25356
rect 46032 25344 46060 25372
rect 46385 25347 46443 25353
rect 46385 25344 46397 25347
rect 35400 25316 37044 25344
rect 46032 25316 46397 25344
rect 35400 25304 35406 25316
rect 27617 25248 27844 25276
rect 27617 25245 27629 25248
rect 27571 25239 27629 25245
rect 24118 25208 24124 25220
rect 23768 25180 24124 25208
rect 22557 25171 22615 25177
rect 24118 25168 24124 25180
rect 24176 25208 24182 25220
rect 25314 25208 25320 25220
rect 24176 25180 25320 25208
rect 24176 25168 24182 25180
rect 25314 25168 25320 25180
rect 25372 25168 25378 25220
rect 22922 25140 22928 25152
rect 22883 25112 22928 25140
rect 22922 25100 22928 25112
rect 22980 25100 22986 25152
rect 27448 25140 27476 25239
rect 27890 25236 27896 25288
rect 27948 25285 27954 25288
rect 27948 25276 27956 25285
rect 29733 25279 29791 25285
rect 27948 25248 27993 25276
rect 27948 25239 27956 25248
rect 29733 25245 29745 25279
rect 29779 25276 29791 25279
rect 31570 25276 31576 25288
rect 29779 25248 30788 25276
rect 31531 25248 31576 25276
rect 29779 25245 29791 25248
rect 29733 25239 29791 25245
rect 27948 25236 27954 25239
rect 27709 25211 27767 25217
rect 27709 25177 27721 25211
rect 27755 25177 27767 25211
rect 27709 25171 27767 25177
rect 27614 25140 27620 25152
rect 27448 25112 27620 25140
rect 27614 25100 27620 25112
rect 27672 25100 27678 25152
rect 27724 25140 27752 25171
rect 27798 25168 27804 25220
rect 27856 25208 27862 25220
rect 27856 25180 27901 25208
rect 27856 25168 27862 25180
rect 29822 25168 29828 25220
rect 29880 25208 29886 25220
rect 29978 25211 30036 25217
rect 29978 25208 29990 25211
rect 29880 25180 29990 25208
rect 29880 25168 29886 25180
rect 29978 25177 29990 25180
rect 30024 25177 30036 25211
rect 30760 25208 30788 25248
rect 31570 25236 31576 25248
rect 31628 25236 31634 25288
rect 35897 25279 35955 25285
rect 35897 25245 35909 25279
rect 35943 25276 35955 25279
rect 36170 25276 36176 25288
rect 35943 25248 36176 25276
rect 35943 25245 35955 25248
rect 35897 25239 35955 25245
rect 36170 25236 36176 25248
rect 36228 25276 36234 25288
rect 36357 25279 36415 25285
rect 36357 25276 36369 25279
rect 36228 25248 36369 25276
rect 36228 25236 36234 25248
rect 36357 25245 36369 25248
rect 36403 25245 36415 25279
rect 36357 25239 36415 25245
rect 36541 25279 36599 25285
rect 36541 25245 36553 25279
rect 36587 25276 36599 25279
rect 36906 25276 36912 25288
rect 36587 25248 36912 25276
rect 36587 25245 36599 25248
rect 36541 25239 36599 25245
rect 36906 25236 36912 25248
rect 36964 25236 36970 25288
rect 37016 25285 37044 25316
rect 46385 25313 46397 25316
rect 46431 25313 46443 25347
rect 46385 25307 46443 25313
rect 37001 25279 37059 25285
rect 37001 25245 37013 25279
rect 37047 25245 37059 25279
rect 37001 25239 37059 25245
rect 37645 25279 37703 25285
rect 37645 25245 37657 25279
rect 37691 25245 37703 25279
rect 39022 25276 39028 25288
rect 38983 25248 39028 25276
rect 37645 25239 37703 25245
rect 31754 25208 31760 25220
rect 30760 25180 31760 25208
rect 29978 25171 30036 25177
rect 31754 25168 31760 25180
rect 31812 25168 31818 25220
rect 35529 25211 35587 25217
rect 35529 25177 35541 25211
rect 35575 25208 35587 25211
rect 35618 25208 35624 25220
rect 35575 25180 35624 25208
rect 35575 25177 35587 25180
rect 35529 25171 35587 25177
rect 35618 25168 35624 25180
rect 35676 25208 35682 25220
rect 36262 25208 36268 25220
rect 35676 25180 36268 25208
rect 35676 25168 35682 25180
rect 36262 25168 36268 25180
rect 36320 25168 36326 25220
rect 36924 25208 36952 25236
rect 37660 25208 37688 25239
rect 39022 25236 39028 25248
rect 39080 25236 39086 25288
rect 41693 25279 41751 25285
rect 41693 25245 41705 25279
rect 41739 25245 41751 25279
rect 42150 25276 42156 25288
rect 42111 25248 42156 25276
rect 41693 25239 41751 25245
rect 38746 25208 38752 25220
rect 36924 25180 37688 25208
rect 38707 25180 38752 25208
rect 38746 25168 38752 25180
rect 38804 25208 38810 25220
rect 41414 25208 41420 25220
rect 38804 25180 41420 25208
rect 38804 25168 38810 25180
rect 41414 25168 41420 25180
rect 41472 25208 41478 25220
rect 41708 25208 41736 25239
rect 42150 25236 42156 25248
rect 42208 25236 42214 25288
rect 42337 25279 42395 25285
rect 42337 25245 42349 25279
rect 42383 25245 42395 25279
rect 45922 25276 45928 25288
rect 45883 25248 45928 25276
rect 42337 25239 42395 25245
rect 41966 25208 41972 25220
rect 41472 25180 41565 25208
rect 41708 25180 41972 25208
rect 41472 25168 41478 25180
rect 41966 25168 41972 25180
rect 42024 25208 42030 25220
rect 42352 25208 42380 25239
rect 45922 25236 45928 25248
rect 45980 25236 45986 25288
rect 46106 25208 46112 25220
rect 42024 25180 42380 25208
rect 46067 25180 46112 25208
rect 42024 25168 42030 25180
rect 46106 25168 46112 25180
rect 46164 25168 46170 25220
rect 28074 25140 28080 25152
rect 27724 25112 28080 25140
rect 28074 25100 28080 25112
rect 28132 25100 28138 25152
rect 30374 25100 30380 25152
rect 30432 25140 30438 25152
rect 31113 25143 31171 25149
rect 31113 25140 31125 25143
rect 30432 25112 31125 25140
rect 30432 25100 30438 25112
rect 31113 25109 31125 25112
rect 31159 25109 31171 25143
rect 31113 25103 31171 25109
rect 31202 25100 31208 25152
rect 31260 25140 31266 25152
rect 31849 25143 31907 25149
rect 31849 25140 31861 25143
rect 31260 25112 31861 25140
rect 31260 25100 31266 25112
rect 31849 25109 31861 25112
rect 31895 25109 31907 25143
rect 37090 25140 37096 25152
rect 37051 25112 37096 25140
rect 31849 25103 31907 25109
rect 37090 25100 37096 25112
rect 37148 25100 37154 25152
rect 37734 25140 37740 25152
rect 37695 25112 37740 25140
rect 37734 25100 37740 25112
rect 37792 25100 37798 25152
rect 38933 25143 38991 25149
rect 38933 25109 38945 25143
rect 38979 25140 38991 25143
rect 39114 25140 39120 25152
rect 38979 25112 39120 25140
rect 38979 25109 38991 25112
rect 38933 25103 38991 25109
rect 39114 25100 39120 25112
rect 39172 25100 39178 25152
rect 41601 25143 41659 25149
rect 41601 25109 41613 25143
rect 41647 25140 41659 25143
rect 42058 25140 42064 25152
rect 41647 25112 42064 25140
rect 41647 25109 41659 25112
rect 41601 25103 41659 25109
rect 42058 25100 42064 25112
rect 42116 25100 42122 25152
rect 42245 25143 42303 25149
rect 42245 25109 42257 25143
rect 42291 25140 42303 25143
rect 42886 25140 42892 25152
rect 42291 25112 42892 25140
rect 42291 25109 42303 25112
rect 42245 25103 42303 25109
rect 42886 25100 42892 25112
rect 42944 25100 42950 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 1762 24896 1768 24948
rect 1820 24936 1826 24948
rect 2409 24939 2467 24945
rect 2409 24936 2421 24939
rect 1820 24908 2421 24936
rect 1820 24896 1826 24908
rect 2409 24905 2421 24908
rect 2455 24905 2467 24939
rect 2409 24899 2467 24905
rect 23661 24939 23719 24945
rect 23661 24905 23673 24939
rect 23707 24936 23719 24939
rect 23842 24936 23848 24948
rect 23707 24908 23848 24936
rect 23707 24905 23719 24908
rect 23661 24899 23719 24905
rect 23842 24896 23848 24908
rect 23900 24896 23906 24948
rect 27890 24896 27896 24948
rect 27948 24936 27954 24948
rect 29822 24936 29828 24948
rect 27948 24908 28994 24936
rect 29783 24908 29828 24936
rect 27948 24896 27954 24908
rect 28966 24868 28994 24908
rect 29822 24896 29828 24908
rect 29880 24896 29886 24948
rect 30926 24896 30932 24948
rect 30984 24936 30990 24948
rect 31113 24939 31171 24945
rect 31113 24936 31125 24939
rect 30984 24908 31125 24936
rect 30984 24896 30990 24908
rect 31113 24905 31125 24908
rect 31159 24905 31171 24939
rect 38746 24936 38752 24948
rect 31113 24899 31171 24905
rect 38672 24908 38752 24936
rect 30742 24868 30748 24880
rect 28966 24840 30748 24868
rect 30742 24828 30748 24840
rect 30800 24828 30806 24880
rect 32490 24828 32496 24880
rect 32548 24868 32554 24880
rect 34790 24868 34796 24880
rect 32548 24840 34796 24868
rect 32548 24828 32554 24840
rect 34790 24828 34796 24840
rect 34848 24868 34854 24880
rect 34848 24840 35848 24868
rect 34848 24828 34854 24840
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24800 2375 24803
rect 2958 24800 2964 24812
rect 2363 24772 2964 24800
rect 2363 24769 2375 24772
rect 2317 24763 2375 24769
rect 2958 24760 2964 24772
rect 3016 24800 3022 24812
rect 3970 24800 3976 24812
rect 3016 24772 3976 24800
rect 3016 24760 3022 24772
rect 3970 24760 3976 24772
rect 4028 24760 4034 24812
rect 22370 24800 22376 24812
rect 22331 24772 22376 24800
rect 22370 24760 22376 24772
rect 22428 24760 22434 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 22738 24800 22744 24812
rect 22603 24772 22744 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 22738 24760 22744 24772
rect 22796 24760 22802 24812
rect 22922 24760 22928 24812
rect 22980 24800 22986 24812
rect 23385 24803 23443 24809
rect 23385 24800 23397 24803
rect 22980 24772 23397 24800
rect 22980 24760 22986 24772
rect 23385 24769 23397 24772
rect 23431 24769 23443 24803
rect 27614 24800 27620 24812
rect 27575 24772 27620 24800
rect 23385 24763 23443 24769
rect 27614 24760 27620 24772
rect 27672 24760 27678 24812
rect 27798 24800 27804 24812
rect 27759 24772 27804 24800
rect 27798 24760 27804 24772
rect 27856 24760 27862 24812
rect 27890 24760 27896 24812
rect 27948 24800 27954 24812
rect 28166 24800 28172 24812
rect 27948 24772 27993 24800
rect 28127 24772 28172 24800
rect 27948 24760 27954 24772
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 30009 24803 30067 24809
rect 30009 24769 30021 24803
rect 30055 24800 30067 24803
rect 30834 24800 30840 24812
rect 30055 24772 30840 24800
rect 30055 24769 30067 24772
rect 30009 24763 30067 24769
rect 30834 24760 30840 24772
rect 30892 24760 30898 24812
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24800 30987 24803
rect 31018 24800 31024 24812
rect 30975 24772 31024 24800
rect 30975 24769 30987 24772
rect 30929 24763 30987 24769
rect 23017 24735 23075 24741
rect 23017 24701 23029 24735
rect 23063 24732 23075 24735
rect 23106 24732 23112 24744
rect 23063 24704 23112 24732
rect 23063 24701 23075 24704
rect 23017 24695 23075 24701
rect 23106 24692 23112 24704
rect 23164 24692 23170 24744
rect 23477 24735 23535 24741
rect 23477 24701 23489 24735
rect 23523 24701 23535 24735
rect 23477 24695 23535 24701
rect 22465 24667 22523 24673
rect 22465 24633 22477 24667
rect 22511 24664 22523 24667
rect 23290 24664 23296 24676
rect 22511 24636 23296 24664
rect 22511 24633 22523 24636
rect 22465 24627 22523 24633
rect 23290 24624 23296 24636
rect 23348 24664 23354 24676
rect 23492 24664 23520 24695
rect 27430 24692 27436 24744
rect 27488 24732 27494 24744
rect 30285 24735 30343 24741
rect 30285 24732 30297 24735
rect 27488 24704 30297 24732
rect 27488 24692 27494 24704
rect 30285 24701 30297 24704
rect 30331 24732 30343 24735
rect 30374 24732 30380 24744
rect 30331 24704 30380 24732
rect 30331 24701 30343 24704
rect 30285 24695 30343 24701
rect 30374 24692 30380 24704
rect 30432 24732 30438 24744
rect 30745 24735 30803 24741
rect 30745 24732 30757 24735
rect 30432 24704 30757 24732
rect 30432 24692 30438 24704
rect 30745 24701 30757 24704
rect 30791 24701 30803 24735
rect 30745 24695 30803 24701
rect 28074 24664 28080 24676
rect 23348 24636 23520 24664
rect 28035 24636 28080 24664
rect 23348 24624 23354 24636
rect 28074 24624 28080 24636
rect 28132 24624 28138 24676
rect 30193 24667 30251 24673
rect 30193 24633 30205 24667
rect 30239 24664 30251 24667
rect 30466 24664 30472 24676
rect 30239 24636 30472 24664
rect 30239 24633 30251 24636
rect 30193 24627 30251 24633
rect 30466 24624 30472 24636
rect 30524 24664 30530 24676
rect 30944 24664 30972 24763
rect 31018 24760 31024 24772
rect 31076 24760 31082 24812
rect 31754 24760 31760 24812
rect 31812 24800 31818 24812
rect 32950 24800 32956 24812
rect 31812 24772 32956 24800
rect 31812 24760 31818 24772
rect 32950 24760 32956 24772
rect 33008 24800 33014 24812
rect 33413 24803 33471 24809
rect 33413 24800 33425 24803
rect 33008 24772 33425 24800
rect 33008 24760 33014 24772
rect 33413 24769 33425 24772
rect 33459 24769 33471 24803
rect 33413 24763 33471 24769
rect 33680 24803 33738 24809
rect 33680 24769 33692 24803
rect 33726 24800 33738 24803
rect 35253 24803 35311 24809
rect 35253 24800 35265 24803
rect 33726 24772 35265 24800
rect 33726 24769 33738 24772
rect 33680 24763 33738 24769
rect 35253 24769 35265 24772
rect 35299 24769 35311 24803
rect 35434 24800 35440 24812
rect 35395 24772 35440 24800
rect 35253 24763 35311 24769
rect 35434 24760 35440 24772
rect 35492 24760 35498 24812
rect 35820 24800 35848 24840
rect 38672 24800 38700 24908
rect 38746 24896 38752 24908
rect 38804 24896 38810 24948
rect 39114 24896 39120 24948
rect 39172 24936 39178 24948
rect 39853 24939 39911 24945
rect 39853 24936 39865 24939
rect 39172 24908 39865 24936
rect 39172 24896 39178 24908
rect 39853 24905 39865 24908
rect 39899 24905 39911 24939
rect 39853 24899 39911 24905
rect 41141 24939 41199 24945
rect 41141 24905 41153 24939
rect 41187 24936 41199 24939
rect 42150 24936 42156 24948
rect 41187 24908 42156 24936
rect 41187 24905 41199 24908
rect 41141 24899 41199 24905
rect 42150 24896 42156 24908
rect 42208 24896 42214 24948
rect 43254 24868 43260 24880
rect 42628 24840 43260 24868
rect 38746 24809 38752 24812
rect 35820 24772 38700 24800
rect 38740 24763 38752 24809
rect 38804 24800 38810 24812
rect 40865 24803 40923 24809
rect 38804 24772 38840 24800
rect 38746 24760 38752 24763
rect 38804 24760 38810 24772
rect 40865 24769 40877 24803
rect 40911 24800 40923 24803
rect 40911 24772 41276 24800
rect 40911 24769 40923 24772
rect 40865 24763 40923 24769
rect 35710 24732 35716 24744
rect 35671 24704 35716 24732
rect 35710 24692 35716 24704
rect 35768 24692 35774 24744
rect 37182 24692 37188 24744
rect 37240 24732 37246 24744
rect 38010 24732 38016 24744
rect 37240 24704 38016 24732
rect 37240 24692 37246 24704
rect 38010 24692 38016 24704
rect 38068 24732 38074 24744
rect 38473 24735 38531 24741
rect 38473 24732 38485 24735
rect 38068 24704 38485 24732
rect 38068 24692 38074 24704
rect 38473 24701 38485 24704
rect 38519 24701 38531 24735
rect 41138 24732 41144 24744
rect 41099 24704 41144 24732
rect 38473 24695 38531 24701
rect 41138 24692 41144 24704
rect 41196 24692 41202 24744
rect 41248 24732 41276 24772
rect 41322 24760 41328 24812
rect 41380 24800 41386 24812
rect 42628 24809 42656 24840
rect 43254 24828 43260 24840
rect 43312 24828 43318 24880
rect 47044 24840 47348 24868
rect 41785 24803 41843 24809
rect 41785 24800 41797 24803
rect 41380 24772 41797 24800
rect 41380 24760 41386 24772
rect 41785 24769 41797 24772
rect 41831 24769 41843 24803
rect 41785 24763 41843 24769
rect 42613 24803 42671 24809
rect 42613 24769 42625 24803
rect 42659 24769 42671 24803
rect 42613 24763 42671 24769
rect 42702 24760 42708 24812
rect 42760 24760 42766 24812
rect 42886 24809 42892 24812
rect 42880 24800 42892 24809
rect 42847 24772 42892 24800
rect 42880 24763 42892 24772
rect 42886 24760 42892 24763
rect 42944 24760 42950 24812
rect 46014 24800 46020 24812
rect 45975 24772 46020 24800
rect 46014 24760 46020 24772
rect 46072 24760 46078 24812
rect 47044 24809 47072 24840
rect 47029 24803 47087 24809
rect 47029 24769 47041 24803
rect 47075 24769 47087 24803
rect 47029 24763 47087 24769
rect 47118 24760 47124 24812
rect 47176 24800 47182 24812
rect 47320 24800 47348 24840
rect 47394 24800 47400 24812
rect 47176 24772 47221 24800
rect 47320 24772 47400 24800
rect 47176 24760 47182 24772
rect 47394 24760 47400 24772
rect 47452 24800 47458 24812
rect 47762 24800 47768 24812
rect 47452 24772 47768 24800
rect 47452 24760 47458 24772
rect 47762 24760 47768 24772
rect 47820 24760 47826 24812
rect 41601 24735 41659 24741
rect 41601 24732 41613 24735
rect 41248 24704 41613 24732
rect 41601 24701 41613 24704
rect 41647 24732 41659 24735
rect 42720 24732 42748 24760
rect 41647 24704 42748 24732
rect 41647 24701 41659 24704
rect 41601 24695 41659 24701
rect 46842 24692 46848 24744
rect 46900 24732 46906 24744
rect 47949 24735 48007 24741
rect 47949 24732 47961 24735
rect 46900 24704 47961 24732
rect 46900 24692 46906 24704
rect 47949 24701 47961 24704
rect 47995 24701 48007 24735
rect 47949 24695 48007 24701
rect 45554 24664 45560 24676
rect 30524 24636 30972 24664
rect 39408 24636 42656 24664
rect 30524 24624 30530 24636
rect 34793 24599 34851 24605
rect 34793 24565 34805 24599
rect 34839 24596 34851 24599
rect 35342 24596 35348 24608
rect 34839 24568 35348 24596
rect 34839 24565 34851 24568
rect 34793 24559 34851 24565
rect 35342 24556 35348 24568
rect 35400 24596 35406 24608
rect 35621 24599 35679 24605
rect 35621 24596 35633 24599
rect 35400 24568 35633 24596
rect 35400 24556 35406 24568
rect 35621 24565 35633 24568
rect 35667 24565 35679 24599
rect 35621 24559 35679 24565
rect 36078 24556 36084 24608
rect 36136 24596 36142 24608
rect 39408 24596 39436 24636
rect 36136 24568 39436 24596
rect 40957 24599 41015 24605
rect 36136 24556 36142 24568
rect 40957 24565 40969 24599
rect 41003 24596 41015 24599
rect 41322 24596 41328 24608
rect 41003 24568 41328 24596
rect 41003 24565 41015 24568
rect 40957 24559 41015 24565
rect 41322 24556 41328 24568
rect 41380 24556 41386 24608
rect 41966 24596 41972 24608
rect 41927 24568 41972 24596
rect 41966 24556 41972 24568
rect 42024 24556 42030 24608
rect 42628 24596 42656 24636
rect 43640 24636 45560 24664
rect 43640 24596 43668 24636
rect 45554 24624 45560 24636
rect 45612 24624 45618 24676
rect 42628 24568 43668 24596
rect 43898 24556 43904 24608
rect 43956 24596 43962 24608
rect 43993 24599 44051 24605
rect 43993 24596 44005 24599
rect 43956 24568 44005 24596
rect 43956 24556 43962 24568
rect 43993 24565 44005 24568
rect 44039 24565 44051 24599
rect 43993 24559 44051 24565
rect 45646 24556 45652 24608
rect 45704 24596 45710 24608
rect 46109 24599 46167 24605
rect 46109 24596 46121 24599
rect 45704 24568 46121 24596
rect 45704 24556 45710 24568
rect 46109 24565 46121 24568
rect 46155 24565 46167 24599
rect 46109 24559 46167 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 24946 24392 24952 24404
rect 24907 24364 24952 24392
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 27798 24352 27804 24404
rect 27856 24392 27862 24404
rect 28813 24395 28871 24401
rect 28813 24392 28825 24395
rect 27856 24364 28825 24392
rect 27856 24352 27862 24364
rect 28813 24361 28825 24364
rect 28859 24361 28871 24395
rect 28813 24355 28871 24361
rect 30009 24395 30067 24401
rect 30009 24361 30021 24395
rect 30055 24392 30067 24395
rect 30374 24392 30380 24404
rect 30055 24364 30380 24392
rect 30055 24361 30067 24364
rect 30009 24355 30067 24361
rect 30374 24352 30380 24364
rect 30432 24352 30438 24404
rect 31570 24392 31576 24404
rect 30484 24364 31576 24392
rect 23290 24256 23296 24268
rect 23251 24228 23296 24256
rect 23290 24216 23296 24228
rect 23348 24216 23354 24268
rect 23661 24259 23719 24265
rect 23661 24225 23673 24259
rect 23707 24256 23719 24259
rect 24964 24256 24992 24352
rect 27706 24284 27712 24336
rect 27764 24284 27770 24336
rect 30484 24324 30512 24364
rect 31570 24352 31576 24364
rect 31628 24392 31634 24404
rect 32033 24395 32091 24401
rect 32033 24392 32045 24395
rect 31628 24364 32045 24392
rect 31628 24352 31634 24364
rect 32033 24361 32045 24364
rect 32079 24361 32091 24395
rect 32033 24355 32091 24361
rect 34885 24395 34943 24401
rect 34885 24361 34897 24395
rect 34931 24392 34943 24395
rect 35434 24392 35440 24404
rect 34931 24364 35440 24392
rect 34931 24361 34943 24364
rect 34885 24355 34943 24361
rect 35434 24352 35440 24364
rect 35492 24352 35498 24404
rect 35710 24352 35716 24404
rect 35768 24392 35774 24404
rect 36725 24395 36783 24401
rect 36725 24392 36737 24395
rect 35768 24364 36737 24392
rect 35768 24352 35774 24364
rect 36725 24361 36737 24364
rect 36771 24392 36783 24395
rect 38657 24395 38715 24401
rect 36771 24364 37872 24392
rect 36771 24361 36783 24364
rect 36725 24355 36783 24361
rect 37734 24324 37740 24336
rect 29840 24296 30512 24324
rect 36648 24296 37740 24324
rect 23707 24228 24992 24256
rect 25041 24259 25099 24265
rect 23707 24225 23719 24228
rect 23661 24219 23719 24225
rect 25041 24225 25053 24259
rect 25087 24256 25099 24259
rect 27724 24256 27752 24284
rect 25087 24228 25728 24256
rect 25087 24225 25099 24228
rect 25041 24219 25099 24225
rect 2038 24148 2044 24200
rect 2096 24188 2102 24200
rect 2317 24191 2375 24197
rect 2317 24188 2329 24191
rect 2096 24160 2329 24188
rect 2096 24148 2102 24160
rect 2317 24157 2329 24160
rect 2363 24157 2375 24191
rect 2317 24151 2375 24157
rect 22186 24148 22192 24200
rect 22244 24188 22250 24200
rect 23014 24188 23020 24200
rect 22244 24160 23020 24188
rect 22244 24148 22250 24160
rect 23014 24148 23020 24160
rect 23072 24188 23078 24200
rect 25700 24197 25728 24228
rect 27172 24228 27752 24256
rect 23753 24191 23811 24197
rect 23753 24188 23765 24191
rect 23072 24160 23765 24188
rect 23072 24148 23078 24160
rect 23753 24157 23765 24160
rect 23799 24188 23811 24191
rect 24765 24191 24823 24197
rect 24765 24188 24777 24191
rect 23799 24160 24777 24188
rect 23799 24157 23811 24160
rect 23753 24151 23811 24157
rect 24765 24157 24777 24160
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 25501 24191 25559 24197
rect 25501 24157 25513 24191
rect 25547 24157 25559 24191
rect 25501 24151 25559 24157
rect 25685 24191 25743 24197
rect 25685 24157 25697 24191
rect 25731 24188 25743 24191
rect 26142 24188 26148 24200
rect 25731 24160 26148 24188
rect 25731 24157 25743 24160
rect 25685 24151 25743 24157
rect 23106 24080 23112 24132
rect 23164 24120 23170 24132
rect 25516 24120 25544 24151
rect 26142 24148 26148 24160
rect 26200 24148 26206 24200
rect 27172 24197 27200 24228
rect 27157 24191 27215 24197
rect 27157 24157 27169 24191
rect 27203 24157 27215 24191
rect 27157 24151 27215 24157
rect 27246 24148 27252 24200
rect 27304 24188 27310 24200
rect 27304 24160 27349 24188
rect 27304 24148 27310 24160
rect 27430 24148 27436 24200
rect 27488 24188 27494 24200
rect 27488 24160 27533 24188
rect 27488 24148 27494 24160
rect 27614 24148 27620 24200
rect 27672 24197 27678 24200
rect 27672 24188 27680 24197
rect 28534 24188 28540 24200
rect 27672 24160 28396 24188
rect 28495 24160 28540 24188
rect 27672 24151 27680 24160
rect 27672 24148 27678 24151
rect 26878 24120 26884 24132
rect 23164 24092 26884 24120
rect 23164 24080 23170 24092
rect 26878 24080 26884 24092
rect 26936 24080 26942 24132
rect 27522 24120 27528 24132
rect 27483 24092 27528 24120
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 28368 24120 28396 24160
rect 28534 24148 28540 24160
rect 28592 24148 28598 24200
rect 28626 24148 28632 24200
rect 28684 24188 28690 24200
rect 28684 24160 28729 24188
rect 28684 24148 28690 24160
rect 29840 24129 29868 24296
rect 32950 24256 32956 24268
rect 32911 24228 32956 24256
rect 32950 24216 32956 24228
rect 33008 24216 33014 24268
rect 30466 24188 30472 24200
rect 30300 24160 30472 24188
rect 29825 24123 29883 24129
rect 29825 24120 29837 24123
rect 28368 24092 29837 24120
rect 29825 24089 29837 24092
rect 29871 24089 29883 24123
rect 29825 24083 29883 24089
rect 30041 24123 30099 24129
rect 30041 24089 30053 24123
rect 30087 24120 30099 24123
rect 30300 24120 30328 24160
rect 30466 24148 30472 24160
rect 30524 24148 30530 24200
rect 30653 24191 30711 24197
rect 30653 24157 30665 24191
rect 30699 24188 30711 24191
rect 31754 24188 31760 24200
rect 30699 24160 31760 24188
rect 30699 24157 30711 24160
rect 30653 24151 30711 24157
rect 31754 24148 31760 24160
rect 31812 24148 31818 24200
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34848 24160 34897 24188
rect 34848 24148 34854 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 35161 24191 35219 24197
rect 35161 24157 35173 24191
rect 35207 24188 35219 24191
rect 35342 24188 35348 24200
rect 35207 24160 35348 24188
rect 35207 24157 35219 24160
rect 35161 24151 35219 24157
rect 35342 24148 35348 24160
rect 35400 24188 35406 24200
rect 36449 24191 36507 24197
rect 36449 24188 36461 24191
rect 35400 24160 36461 24188
rect 35400 24148 35406 24160
rect 36449 24157 36461 24160
rect 36495 24157 36507 24191
rect 36449 24151 36507 24157
rect 36541 24191 36599 24197
rect 36541 24157 36553 24191
rect 36587 24188 36599 24191
rect 36648 24188 36676 24296
rect 37734 24284 37740 24296
rect 37792 24284 37798 24336
rect 37844 24256 37872 24364
rect 38657 24361 38669 24395
rect 38703 24392 38715 24395
rect 38746 24392 38752 24404
rect 38703 24364 38752 24392
rect 38703 24361 38715 24364
rect 38657 24355 38715 24361
rect 38746 24352 38752 24364
rect 38804 24352 38810 24404
rect 41966 24352 41972 24404
rect 42024 24392 42030 24404
rect 42429 24395 42487 24401
rect 42429 24392 42441 24395
rect 42024 24364 42441 24392
rect 42024 24352 42030 24364
rect 42429 24361 42441 24364
rect 42475 24361 42487 24395
rect 44174 24392 44180 24404
rect 42429 24355 42487 24361
rect 42536 24364 44180 24392
rect 37918 24284 37924 24336
rect 37976 24324 37982 24336
rect 41138 24324 41144 24336
rect 37976 24296 41144 24324
rect 37976 24284 37982 24296
rect 41138 24284 41144 24296
rect 41196 24284 41202 24336
rect 37476 24228 37872 24256
rect 36587 24160 36676 24188
rect 36817 24191 36875 24197
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 36817 24157 36829 24191
rect 36863 24188 36875 24191
rect 37090 24188 37096 24200
rect 36863 24160 37096 24188
rect 36863 24157 36875 24160
rect 36817 24151 36875 24157
rect 30087 24092 30328 24120
rect 30087 24089 30099 24092
rect 30041 24083 30099 24089
rect 30374 24080 30380 24132
rect 30432 24120 30438 24132
rect 30898 24123 30956 24129
rect 30898 24120 30910 24123
rect 30432 24092 30910 24120
rect 30432 24080 30438 24092
rect 30898 24089 30910 24092
rect 30944 24089 30956 24123
rect 30898 24083 30956 24089
rect 33220 24123 33278 24129
rect 33220 24089 33232 24123
rect 33266 24120 33278 24123
rect 33778 24120 33784 24132
rect 33266 24092 33784 24120
rect 33266 24089 33278 24092
rect 33220 24083 33278 24089
rect 33778 24080 33784 24092
rect 33836 24080 33842 24132
rect 35986 24080 35992 24132
rect 36044 24120 36050 24132
rect 36556 24120 36584 24151
rect 37090 24148 37096 24160
rect 37148 24148 37154 24200
rect 37476 24197 37504 24228
rect 38654 24216 38660 24268
rect 38712 24256 38718 24268
rect 39022 24256 39028 24268
rect 38712 24228 39028 24256
rect 38712 24216 38718 24228
rect 39022 24216 39028 24228
rect 39080 24256 39086 24268
rect 40126 24256 40132 24268
rect 39080 24228 40132 24256
rect 39080 24216 39086 24228
rect 40126 24216 40132 24228
rect 40184 24216 40190 24268
rect 42058 24216 42064 24268
rect 42116 24256 42122 24268
rect 42536 24265 42564 24364
rect 44174 24352 44180 24364
rect 44232 24392 44238 24404
rect 44637 24395 44695 24401
rect 44637 24392 44649 24395
rect 44232 24364 44649 24392
rect 44232 24352 44238 24364
rect 44637 24361 44649 24364
rect 44683 24361 44695 24395
rect 44637 24355 44695 24361
rect 45925 24395 45983 24401
rect 45925 24361 45937 24395
rect 45971 24392 45983 24395
rect 46106 24392 46112 24404
rect 45971 24364 46112 24392
rect 45971 24361 45983 24364
rect 45925 24355 45983 24361
rect 46106 24352 46112 24364
rect 46164 24352 46170 24404
rect 42521 24259 42579 24265
rect 42521 24256 42533 24259
rect 42116 24228 42533 24256
rect 42116 24216 42122 24228
rect 42521 24225 42533 24228
rect 42567 24225 42579 24259
rect 43254 24256 43260 24268
rect 43215 24228 43260 24256
rect 42521 24219 42579 24225
rect 43254 24216 43260 24228
rect 43312 24216 43318 24268
rect 37461 24191 37519 24197
rect 37461 24157 37473 24191
rect 37507 24157 37519 24191
rect 37461 24151 37519 24157
rect 37553 24191 37611 24197
rect 37553 24157 37565 24191
rect 37599 24157 37611 24191
rect 37734 24188 37740 24200
rect 37695 24160 37740 24188
rect 37553 24151 37611 24157
rect 36044 24092 36584 24120
rect 37108 24120 37136 24148
rect 37568 24120 37596 24151
rect 37734 24148 37740 24160
rect 37792 24148 37798 24200
rect 37829 24191 37887 24197
rect 37829 24157 37841 24191
rect 37875 24157 37887 24191
rect 38838 24188 38844 24200
rect 38799 24160 38844 24188
rect 37829 24151 37887 24157
rect 37108 24092 37596 24120
rect 36044 24080 36050 24092
rect 23934 24052 23940 24064
rect 23895 24024 23940 24052
rect 23934 24012 23940 24024
rect 23992 24012 23998 24064
rect 24578 24052 24584 24064
rect 24539 24024 24584 24052
rect 24578 24012 24584 24024
rect 24636 24012 24642 24064
rect 25498 24012 25504 24064
rect 25556 24052 25562 24064
rect 25593 24055 25651 24061
rect 25593 24052 25605 24055
rect 25556 24024 25605 24052
rect 25556 24012 25562 24024
rect 25593 24021 25605 24024
rect 25639 24021 25651 24055
rect 27798 24052 27804 24064
rect 27759 24024 27804 24052
rect 25593 24015 25651 24021
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 30193 24055 30251 24061
rect 30193 24021 30205 24055
rect 30239 24052 30251 24055
rect 30466 24052 30472 24064
rect 30239 24024 30472 24052
rect 30239 24021 30251 24024
rect 30193 24015 30251 24021
rect 30466 24012 30472 24024
rect 30524 24012 30530 24064
rect 34333 24055 34391 24061
rect 34333 24021 34345 24055
rect 34379 24052 34391 24055
rect 34606 24052 34612 24064
rect 34379 24024 34612 24052
rect 34379 24021 34391 24024
rect 34333 24015 34391 24021
rect 34606 24012 34612 24024
rect 34664 24052 34670 24064
rect 35069 24055 35127 24061
rect 35069 24052 35081 24055
rect 34664 24024 35081 24052
rect 34664 24012 34670 24024
rect 35069 24021 35081 24024
rect 35115 24052 35127 24055
rect 35710 24052 35716 24064
rect 35115 24024 35716 24052
rect 35115 24021 35127 24024
rect 35069 24015 35127 24021
rect 35710 24012 35716 24024
rect 35768 24012 35774 24064
rect 36265 24055 36323 24061
rect 36265 24021 36277 24055
rect 36311 24052 36323 24055
rect 36906 24052 36912 24064
rect 36311 24024 36912 24052
rect 36311 24021 36323 24024
rect 36265 24015 36323 24021
rect 36906 24012 36912 24024
rect 36964 24012 36970 24064
rect 37274 24052 37280 24064
rect 37235 24024 37280 24052
rect 37274 24012 37280 24024
rect 37332 24012 37338 24064
rect 37844 24052 37872 24151
rect 38838 24148 38844 24160
rect 38896 24148 38902 24200
rect 39114 24188 39120 24200
rect 39075 24160 39120 24188
rect 39114 24148 39120 24160
rect 39172 24148 39178 24200
rect 42242 24188 42248 24200
rect 42203 24160 42248 24188
rect 42242 24148 42248 24160
rect 42300 24148 42306 24200
rect 45646 24148 45652 24200
rect 45704 24188 45710 24200
rect 45833 24191 45891 24197
rect 45833 24188 45845 24191
rect 45704 24160 45845 24188
rect 45704 24148 45710 24160
rect 45833 24157 45845 24160
rect 45879 24188 45891 24191
rect 46658 24188 46664 24200
rect 45879 24160 46664 24188
rect 45879 24157 45891 24160
rect 45833 24151 45891 24157
rect 46658 24148 46664 24160
rect 46716 24148 46722 24200
rect 42061 24123 42119 24129
rect 42061 24089 42073 24123
rect 42107 24120 42119 24123
rect 43502 24123 43560 24129
rect 43502 24120 43514 24123
rect 42107 24092 43514 24120
rect 42107 24089 42119 24092
rect 42061 24083 42119 24089
rect 43502 24089 43514 24092
rect 43548 24089 43560 24123
rect 43502 24083 43560 24089
rect 41138 24052 41144 24064
rect 37844 24024 41144 24052
rect 41138 24012 41144 24024
rect 41196 24012 41202 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 26237 23851 26295 23857
rect 26237 23848 26249 23851
rect 22296 23820 26249 23848
rect 3510 23740 3516 23792
rect 3568 23780 3574 23792
rect 3568 23752 6914 23780
rect 3568 23740 3574 23752
rect 2038 23712 2044 23724
rect 1999 23684 2044 23712
rect 2038 23672 2044 23684
rect 2096 23672 2102 23724
rect 2222 23644 2228 23656
rect 2183 23616 2228 23644
rect 2222 23604 2228 23616
rect 2280 23604 2286 23656
rect 2774 23644 2780 23656
rect 2735 23616 2780 23644
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 6886 23576 6914 23752
rect 22296 23721 22324 23820
rect 26237 23817 26249 23820
rect 26283 23848 26295 23851
rect 27246 23848 27252 23860
rect 26283 23820 27252 23848
rect 26283 23817 26295 23820
rect 26237 23811 26295 23817
rect 27246 23808 27252 23820
rect 27304 23848 27310 23860
rect 27982 23848 27988 23860
rect 27304 23820 27988 23848
rect 27304 23808 27310 23820
rect 27982 23808 27988 23820
rect 28040 23808 28046 23860
rect 30374 23848 30380 23860
rect 30335 23820 30380 23848
rect 30374 23808 30380 23820
rect 30432 23808 30438 23860
rect 30558 23808 30564 23860
rect 30616 23848 30622 23860
rect 31129 23851 31187 23857
rect 31129 23848 31141 23851
rect 30616 23820 31141 23848
rect 30616 23808 30622 23820
rect 31129 23817 31141 23820
rect 31175 23817 31187 23851
rect 31294 23848 31300 23860
rect 31255 23820 31300 23848
rect 31129 23811 31187 23817
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 33778 23848 33784 23860
rect 33739 23820 33784 23848
rect 33778 23808 33784 23820
rect 33836 23808 33842 23860
rect 37734 23808 37740 23860
rect 37792 23848 37798 23860
rect 38933 23851 38991 23857
rect 38933 23848 38945 23851
rect 37792 23820 38945 23848
rect 37792 23808 37798 23820
rect 38933 23817 38945 23820
rect 38979 23817 38991 23851
rect 38933 23811 38991 23817
rect 40126 23808 40132 23860
rect 40184 23857 40190 23860
rect 40184 23851 40203 23857
rect 40191 23817 40203 23851
rect 40184 23811 40203 23817
rect 40313 23851 40371 23857
rect 40313 23817 40325 23851
rect 40359 23848 40371 23851
rect 40770 23848 40776 23860
rect 40359 23820 40776 23848
rect 40359 23817 40371 23820
rect 40313 23811 40371 23817
rect 40184 23808 40190 23811
rect 40770 23808 40776 23820
rect 40828 23848 40834 23860
rect 41322 23848 41328 23860
rect 40828 23820 41328 23848
rect 40828 23808 40834 23820
rect 41322 23808 41328 23820
rect 41380 23808 41386 23860
rect 22738 23740 22744 23792
rect 22796 23780 22802 23792
rect 22796 23752 23520 23780
rect 22796 23740 22802 23752
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 22370 23672 22376 23724
rect 22428 23712 22434 23724
rect 23492 23721 23520 23752
rect 30742 23740 30748 23792
rect 30800 23780 30806 23792
rect 30926 23780 30932 23792
rect 30800 23752 30932 23780
rect 30800 23740 30806 23752
rect 30926 23740 30932 23752
rect 30984 23740 30990 23792
rect 35342 23740 35348 23792
rect 35400 23780 35406 23792
rect 36173 23783 36231 23789
rect 36173 23780 36185 23783
rect 35400 23752 36185 23780
rect 35400 23740 35406 23752
rect 36173 23749 36185 23752
rect 36219 23749 36231 23783
rect 39942 23780 39948 23792
rect 39903 23752 39948 23780
rect 36173 23743 36231 23749
rect 39942 23740 39948 23752
rect 40000 23740 40006 23792
rect 41785 23783 41843 23789
rect 41785 23749 41797 23783
rect 41831 23780 41843 23783
rect 44082 23780 44088 23792
rect 41831 23752 44088 23780
rect 41831 23749 41843 23752
rect 41785 23743 41843 23749
rect 44082 23740 44088 23752
rect 44140 23740 44146 23792
rect 47213 23783 47271 23789
rect 47213 23749 47225 23783
rect 47259 23780 47271 23783
rect 48038 23780 48044 23792
rect 47259 23752 48044 23780
rect 47259 23749 47271 23752
rect 47213 23743 47271 23749
rect 48038 23740 48044 23752
rect 48096 23740 48102 23792
rect 23385 23715 23443 23721
rect 23385 23712 23397 23715
rect 22428 23684 23397 23712
rect 22428 23672 22434 23684
rect 23385 23681 23397 23684
rect 23431 23681 23443 23715
rect 23385 23675 23443 23681
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23681 23535 23715
rect 23477 23675 23535 23681
rect 23569 23715 23627 23721
rect 23569 23681 23581 23715
rect 23615 23712 23627 23715
rect 24578 23712 24584 23724
rect 23615 23684 24584 23712
rect 23615 23681 23627 23684
rect 23569 23675 23627 23681
rect 24578 23672 24584 23684
rect 24636 23672 24642 23724
rect 24854 23672 24860 23724
rect 24912 23712 24918 23724
rect 25225 23715 25283 23721
rect 25225 23712 25237 23715
rect 24912 23684 25237 23712
rect 24912 23672 24918 23684
rect 25225 23681 25237 23684
rect 25271 23681 25283 23715
rect 25225 23675 25283 23681
rect 25314 23672 25320 23724
rect 25372 23712 25378 23724
rect 25498 23712 25504 23724
rect 25372 23684 25417 23712
rect 25459 23684 25504 23712
rect 25372 23672 25378 23684
rect 25498 23672 25504 23684
rect 25556 23672 25562 23724
rect 26142 23712 26148 23724
rect 26103 23684 26148 23712
rect 26142 23672 26148 23684
rect 26200 23672 26206 23724
rect 30285 23715 30343 23721
rect 30285 23681 30297 23715
rect 30331 23681 30343 23715
rect 30466 23712 30472 23724
rect 30427 23684 30472 23712
rect 30285 23675 30343 23681
rect 22186 23644 22192 23656
rect 22147 23616 22192 23644
rect 22186 23604 22192 23616
rect 22244 23604 22250 23656
rect 23198 23644 23204 23656
rect 22664 23616 23204 23644
rect 22664 23585 22692 23616
rect 23198 23604 23204 23616
rect 23256 23644 23262 23656
rect 23293 23647 23351 23653
rect 23293 23644 23305 23647
rect 23256 23616 23305 23644
rect 23256 23604 23262 23616
rect 23293 23613 23305 23616
rect 23339 23613 23351 23647
rect 23293 23607 23351 23613
rect 25593 23647 25651 23653
rect 25593 23613 25605 23647
rect 25639 23644 25651 23647
rect 26970 23644 26976 23656
rect 25639 23616 26976 23644
rect 25639 23613 25651 23616
rect 25593 23607 25651 23613
rect 26970 23604 26976 23616
rect 27028 23604 27034 23656
rect 27706 23644 27712 23656
rect 27667 23616 27712 23644
rect 27706 23604 27712 23616
rect 27764 23604 27770 23656
rect 27893 23647 27951 23653
rect 27893 23613 27905 23647
rect 27939 23644 27951 23647
rect 28442 23644 28448 23656
rect 27939 23616 28448 23644
rect 27939 23613 27951 23616
rect 27893 23607 27951 23613
rect 28442 23604 28448 23616
rect 28500 23604 28506 23656
rect 28537 23647 28595 23653
rect 28537 23613 28549 23647
rect 28583 23613 28595 23647
rect 30300 23644 30328 23675
rect 30466 23672 30472 23684
rect 30524 23672 30530 23724
rect 33686 23712 33692 23724
rect 33647 23684 33692 23712
rect 33686 23672 33692 23684
rect 33744 23672 33750 23724
rect 33873 23715 33931 23721
rect 33873 23681 33885 23715
rect 33919 23712 33931 23715
rect 34606 23712 34612 23724
rect 33919 23684 34612 23712
rect 33919 23681 33931 23684
rect 33873 23675 33931 23681
rect 34606 23672 34612 23684
rect 34664 23672 34670 23724
rect 35986 23712 35992 23724
rect 35947 23684 35992 23712
rect 35986 23672 35992 23684
rect 36044 23672 36050 23724
rect 36262 23712 36268 23724
rect 36223 23684 36268 23712
rect 36262 23672 36268 23684
rect 36320 23672 36326 23724
rect 36354 23672 36360 23724
rect 36412 23712 36418 23724
rect 37461 23715 37519 23721
rect 36412 23684 36457 23712
rect 36412 23672 36418 23684
rect 37461 23681 37473 23715
rect 37507 23712 37519 23715
rect 37642 23712 37648 23724
rect 37507 23684 37648 23712
rect 37507 23681 37519 23684
rect 37461 23675 37519 23681
rect 37642 23672 37648 23684
rect 37700 23672 37706 23724
rect 38841 23715 38899 23721
rect 38841 23681 38853 23715
rect 38887 23681 38899 23715
rect 38841 23675 38899 23681
rect 31202 23644 31208 23656
rect 30300 23616 31208 23644
rect 28537 23607 28595 23613
rect 22649 23579 22707 23585
rect 6886 23548 22094 23576
rect 22066 23508 22094 23548
rect 22649 23545 22661 23579
rect 22695 23545 22707 23579
rect 28552 23576 28580 23607
rect 31202 23604 31208 23616
rect 31260 23604 31266 23656
rect 37737 23647 37795 23653
rect 37737 23613 37749 23647
rect 37783 23644 37795 23647
rect 37918 23644 37924 23656
rect 37783 23616 37924 23644
rect 37783 23613 37795 23616
rect 37737 23607 37795 23613
rect 37918 23604 37924 23616
rect 37976 23604 37982 23656
rect 38856 23644 38884 23675
rect 40034 23672 40040 23724
rect 40092 23712 40098 23724
rect 41417 23715 41475 23721
rect 41417 23712 41429 23715
rect 40092 23684 41429 23712
rect 40092 23672 40098 23684
rect 41417 23681 41429 23684
rect 41463 23681 41475 23715
rect 41417 23675 41475 23681
rect 41506 23672 41512 23724
rect 41564 23712 41570 23724
rect 41564 23684 41609 23712
rect 41564 23672 41570 23684
rect 41690 23672 41696 23724
rect 41748 23712 41754 23724
rect 41923 23715 41981 23721
rect 41748 23684 41793 23712
rect 41748 23672 41754 23684
rect 41923 23681 41935 23715
rect 41969 23712 41981 23715
rect 42794 23712 42800 23724
rect 41969 23684 42800 23712
rect 41969 23681 41981 23684
rect 41923 23675 41981 23681
rect 42794 23672 42800 23684
rect 42852 23712 42858 23724
rect 43898 23712 43904 23724
rect 42852 23684 43904 23712
rect 42852 23672 42858 23684
rect 43898 23672 43904 23684
rect 43956 23672 43962 23724
rect 42058 23644 42064 23656
rect 38856 23616 42064 23644
rect 42058 23604 42064 23616
rect 42116 23604 42122 23656
rect 45370 23644 45376 23656
rect 45331 23616 45376 23644
rect 45370 23604 45376 23616
rect 45428 23604 45434 23656
rect 45554 23644 45560 23656
rect 45515 23616 45560 23644
rect 45554 23604 45560 23616
rect 45612 23604 45618 23656
rect 22649 23539 22707 23545
rect 22756 23548 28580 23576
rect 22756 23508 22784 23548
rect 39482 23536 39488 23588
rect 39540 23576 39546 23588
rect 41506 23576 41512 23588
rect 39540 23548 41512 23576
rect 39540 23536 39546 23548
rect 41506 23536 41512 23548
rect 41564 23576 41570 23588
rect 41966 23576 41972 23588
rect 41564 23548 41972 23576
rect 41564 23536 41570 23548
rect 41966 23536 41972 23548
rect 42024 23536 42030 23588
rect 23106 23508 23112 23520
rect 22066 23480 22784 23508
rect 23067 23480 23112 23508
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25593 23511 25651 23517
rect 25593 23508 25605 23511
rect 25004 23480 25605 23508
rect 25004 23468 25010 23480
rect 25593 23477 25605 23480
rect 25639 23477 25651 23511
rect 25593 23471 25651 23477
rect 28074 23468 28080 23520
rect 28132 23508 28138 23520
rect 31113 23511 31171 23517
rect 31113 23508 31125 23511
rect 28132 23480 31125 23508
rect 28132 23468 28138 23480
rect 31113 23477 31125 23480
rect 31159 23508 31171 23511
rect 31386 23508 31392 23520
rect 31159 23480 31392 23508
rect 31159 23477 31171 23480
rect 31113 23471 31171 23477
rect 31386 23468 31392 23480
rect 31444 23468 31450 23520
rect 36541 23511 36599 23517
rect 36541 23477 36553 23511
rect 36587 23508 36599 23511
rect 36630 23508 36636 23520
rect 36587 23480 36636 23508
rect 36587 23477 36599 23480
rect 36541 23471 36599 23477
rect 36630 23468 36636 23480
rect 36688 23468 36694 23520
rect 37550 23508 37556 23520
rect 37511 23480 37556 23508
rect 37550 23468 37556 23480
rect 37608 23468 37614 23520
rect 37645 23511 37703 23517
rect 37645 23477 37657 23511
rect 37691 23508 37703 23511
rect 38286 23508 38292 23520
rect 37691 23480 38292 23508
rect 37691 23477 37703 23480
rect 37645 23471 37703 23477
rect 38286 23468 38292 23480
rect 38344 23468 38350 23520
rect 39114 23468 39120 23520
rect 39172 23508 39178 23520
rect 40129 23511 40187 23517
rect 40129 23508 40141 23511
rect 39172 23480 40141 23508
rect 39172 23468 39178 23480
rect 40129 23477 40141 23480
rect 40175 23508 40187 23511
rect 40218 23508 40224 23520
rect 40175 23480 40224 23508
rect 40175 23477 40187 23480
rect 40129 23471 40187 23477
rect 40218 23468 40224 23480
rect 40276 23468 40282 23520
rect 42061 23511 42119 23517
rect 42061 23477 42073 23511
rect 42107 23508 42119 23511
rect 43806 23508 43812 23520
rect 42107 23480 43812 23508
rect 42107 23477 42119 23480
rect 42061 23471 42119 23477
rect 43806 23468 43812 23480
rect 43864 23468 43870 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 2222 23264 2228 23316
rect 2280 23304 2286 23316
rect 2501 23307 2559 23313
rect 2501 23304 2513 23307
rect 2280 23276 2513 23304
rect 2280 23264 2286 23276
rect 2501 23273 2513 23276
rect 2547 23273 2559 23307
rect 2501 23267 2559 23273
rect 23477 23307 23535 23313
rect 23477 23273 23489 23307
rect 23523 23304 23535 23307
rect 24854 23304 24860 23316
rect 23523 23276 24860 23304
rect 23523 23273 23535 23276
rect 23477 23267 23535 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 26053 23307 26111 23313
rect 26053 23273 26065 23307
rect 26099 23304 26111 23307
rect 26142 23304 26148 23316
rect 26099 23276 26148 23304
rect 26099 23273 26111 23276
rect 26053 23267 26111 23273
rect 26142 23264 26148 23276
rect 26200 23264 26206 23316
rect 27890 23264 27896 23316
rect 27948 23304 27954 23316
rect 27985 23307 28043 23313
rect 27985 23304 27997 23307
rect 27948 23276 27997 23304
rect 27948 23264 27954 23276
rect 27985 23273 27997 23276
rect 28031 23273 28043 23307
rect 28534 23304 28540 23316
rect 28495 23276 28540 23304
rect 27985 23267 28043 23273
rect 28534 23264 28540 23276
rect 28592 23264 28598 23316
rect 34698 23264 34704 23316
rect 34756 23304 34762 23316
rect 35069 23307 35127 23313
rect 35069 23304 35081 23307
rect 34756 23276 35081 23304
rect 34756 23264 34762 23276
rect 35069 23273 35081 23276
rect 35115 23273 35127 23307
rect 35069 23267 35127 23273
rect 45554 23264 45560 23316
rect 45612 23304 45618 23316
rect 45741 23307 45799 23313
rect 45741 23304 45753 23307
rect 45612 23276 45753 23304
rect 45612 23264 45618 23276
rect 45741 23273 45753 23276
rect 45787 23273 45799 23307
rect 45741 23267 45799 23273
rect 27798 23236 27804 23248
rect 27356 23208 27804 23236
rect 23293 23171 23351 23177
rect 23293 23137 23305 23171
rect 23339 23168 23351 23171
rect 23934 23168 23940 23180
rect 23339 23140 23940 23168
rect 23339 23137 23351 23140
rect 23293 23131 23351 23137
rect 23934 23128 23940 23140
rect 23992 23128 23998 23180
rect 2406 23100 2412 23112
rect 2367 23072 2412 23100
rect 2406 23060 2412 23072
rect 2464 23060 2470 23112
rect 23198 23100 23204 23112
rect 23159 23072 23204 23100
rect 23198 23060 23204 23072
rect 23256 23060 23262 23112
rect 24394 23060 24400 23112
rect 24452 23100 24458 23112
rect 24946 23109 24952 23112
rect 24673 23103 24731 23109
rect 24673 23100 24685 23103
rect 24452 23072 24685 23100
rect 24452 23060 24458 23072
rect 24673 23069 24685 23072
rect 24719 23069 24731 23103
rect 24940 23100 24952 23109
rect 24907 23072 24952 23100
rect 24673 23063 24731 23069
rect 24940 23063 24952 23072
rect 24946 23060 24952 23063
rect 25004 23060 25010 23112
rect 26970 23100 26976 23112
rect 26931 23072 26976 23100
rect 26970 23060 26976 23072
rect 27028 23060 27034 23112
rect 27062 23060 27068 23112
rect 27120 23100 27126 23112
rect 27249 23103 27307 23109
rect 27120 23072 27165 23100
rect 27120 23060 27126 23072
rect 27249 23069 27261 23103
rect 27295 23100 27307 23103
rect 27356 23100 27384 23208
rect 27798 23196 27804 23208
rect 27856 23196 27862 23248
rect 30558 23236 30564 23248
rect 28644 23208 30564 23236
rect 28644 23180 28672 23208
rect 30558 23196 30564 23208
rect 30616 23196 30622 23248
rect 31294 23236 31300 23248
rect 30668 23208 31300 23236
rect 27525 23171 27583 23177
rect 27525 23137 27537 23171
rect 27571 23168 27583 23171
rect 27706 23168 27712 23180
rect 27571 23140 27712 23168
rect 27571 23137 27583 23140
rect 27525 23131 27583 23137
rect 27706 23128 27712 23140
rect 27764 23128 27770 23180
rect 28626 23168 28632 23180
rect 28587 23140 28632 23168
rect 28626 23128 28632 23140
rect 28684 23128 28690 23180
rect 30668 23168 30696 23208
rect 31294 23196 31300 23208
rect 31352 23196 31358 23248
rect 34790 23196 34796 23248
rect 34848 23236 34854 23248
rect 35253 23239 35311 23245
rect 35253 23236 35265 23239
rect 34848 23208 35265 23236
rect 34848 23196 34854 23208
rect 35253 23205 35265 23208
rect 35299 23236 35311 23239
rect 37642 23236 37648 23248
rect 35299 23208 37648 23236
rect 35299 23205 35311 23208
rect 35253 23199 35311 23205
rect 37642 23196 37648 23208
rect 37700 23196 37706 23248
rect 40037 23239 40095 23245
rect 40037 23205 40049 23239
rect 40083 23236 40095 23239
rect 40865 23239 40923 23245
rect 40865 23236 40877 23239
rect 40083 23208 40877 23236
rect 40083 23205 40095 23208
rect 40037 23199 40095 23205
rect 40865 23205 40877 23208
rect 40911 23205 40923 23239
rect 40865 23199 40923 23205
rect 30576 23140 30696 23168
rect 30837 23171 30895 23177
rect 27295 23072 27384 23100
rect 27433 23103 27491 23109
rect 27295 23069 27307 23072
rect 27249 23063 27307 23069
rect 27433 23069 27445 23103
rect 27479 23100 27491 23103
rect 27798 23100 27804 23112
rect 27479 23072 27804 23100
rect 27479 23069 27491 23072
rect 27433 23063 27491 23069
rect 27798 23060 27804 23072
rect 27856 23060 27862 23112
rect 28166 23100 28172 23112
rect 27908 23072 28172 23100
rect 27341 23035 27399 23041
rect 27341 23001 27353 23035
rect 27387 23032 27399 23035
rect 27908 23032 27936 23072
rect 28166 23060 28172 23072
rect 28224 23060 28230 23112
rect 30576 23109 30604 23140
rect 30837 23137 30849 23171
rect 30883 23168 30895 23171
rect 36449 23171 36507 23177
rect 30883 23140 31432 23168
rect 30883 23137 30895 23140
rect 30837 23131 30895 23137
rect 30561 23103 30619 23109
rect 30561 23069 30573 23103
rect 30607 23069 30619 23103
rect 30561 23063 30619 23069
rect 30650 23060 30656 23112
rect 30708 23100 30714 23112
rect 31294 23100 31300 23112
rect 30708 23072 30753 23100
rect 31255 23072 31300 23100
rect 30708 23060 30714 23072
rect 31294 23060 31300 23072
rect 31352 23060 31358 23112
rect 31404 23100 31432 23140
rect 36449 23137 36461 23171
rect 36495 23168 36507 23171
rect 41690 23168 41696 23180
rect 36495 23140 37872 23168
rect 36495 23137 36507 23140
rect 36449 23131 36507 23137
rect 33686 23100 33692 23112
rect 31404 23072 33692 23100
rect 33686 23060 33692 23072
rect 33744 23100 33750 23112
rect 33962 23100 33968 23112
rect 33744 23072 33968 23100
rect 33744 23060 33750 23072
rect 33962 23060 33968 23072
rect 34020 23060 34026 23112
rect 36630 23100 36636 23112
rect 36591 23072 36636 23100
rect 36630 23060 36636 23072
rect 36688 23060 36694 23112
rect 36906 23100 36912 23112
rect 36867 23072 36912 23100
rect 36906 23060 36912 23072
rect 36964 23060 36970 23112
rect 37550 23100 37556 23112
rect 37511 23072 37556 23100
rect 37550 23060 37556 23072
rect 37608 23060 37614 23112
rect 37844 23109 37872 23140
rect 40052 23140 41696 23168
rect 37829 23103 37887 23109
rect 37829 23069 37841 23103
rect 37875 23069 37887 23103
rect 38286 23100 38292 23112
rect 38247 23072 38292 23100
rect 37829 23063 37887 23069
rect 38286 23060 38292 23072
rect 38344 23060 38350 23112
rect 38470 23100 38476 23112
rect 38431 23072 38476 23100
rect 38470 23060 38476 23072
rect 38528 23060 38534 23112
rect 31542 23035 31600 23041
rect 31542 23032 31554 23035
rect 27387 23004 27936 23032
rect 31036 23004 31554 23032
rect 27387 23001 27399 23004
rect 27341 22995 27399 23001
rect 27798 22924 27804 22976
rect 27856 22964 27862 22976
rect 28169 22967 28227 22973
rect 28169 22964 28181 22967
rect 27856 22936 28181 22964
rect 27856 22924 27862 22936
rect 28169 22933 28181 22936
rect 28215 22964 28227 22967
rect 29914 22964 29920 22976
rect 28215 22936 29920 22964
rect 28215 22933 28227 22936
rect 28169 22927 28227 22933
rect 29914 22924 29920 22936
rect 29972 22924 29978 22976
rect 30561 22967 30619 22973
rect 30561 22933 30573 22967
rect 30607 22964 30619 22967
rect 31036 22964 31064 23004
rect 31542 23001 31554 23004
rect 31588 23001 31600 23035
rect 31542 22995 31600 23001
rect 34606 22992 34612 23044
rect 34664 23032 34670 23044
rect 34885 23035 34943 23041
rect 34885 23032 34897 23035
rect 34664 23004 34897 23032
rect 34664 22992 34670 23004
rect 34885 23001 34897 23004
rect 34931 23001 34943 23035
rect 34885 22995 34943 23001
rect 35101 23035 35159 23041
rect 35101 23001 35113 23035
rect 35147 23032 35159 23035
rect 35342 23032 35348 23044
rect 35147 23004 35348 23032
rect 35147 23001 35159 23004
rect 35101 22995 35159 23001
rect 35342 22992 35348 23004
rect 35400 22992 35406 23044
rect 36817 23035 36875 23041
rect 36817 23001 36829 23035
rect 36863 23032 36875 23035
rect 37274 23032 37280 23044
rect 36863 23004 37280 23032
rect 36863 23001 36875 23004
rect 36817 22995 36875 23001
rect 37274 22992 37280 23004
rect 37332 22992 37338 23044
rect 39298 22992 39304 23044
rect 39356 23032 39362 23044
rect 39942 23032 39948 23044
rect 39356 23004 39948 23032
rect 39356 22992 39362 23004
rect 39942 22992 39948 23004
rect 40000 23032 40006 23044
rect 40052 23041 40080 23140
rect 41690 23128 41696 23140
rect 41748 23128 41754 23180
rect 42702 23128 42708 23180
rect 42760 23168 42766 23180
rect 43254 23168 43260 23180
rect 42760 23140 43260 23168
rect 42760 23128 42766 23140
rect 43254 23128 43260 23140
rect 43312 23128 43318 23180
rect 44082 23168 44088 23180
rect 44043 23140 44088 23168
rect 44082 23128 44088 23140
rect 44140 23128 44146 23180
rect 44174 23128 44180 23180
rect 44232 23168 44238 23180
rect 44232 23140 44277 23168
rect 44232 23128 44238 23140
rect 40126 23060 40132 23112
rect 40184 23100 40190 23112
rect 40313 23103 40371 23109
rect 40313 23100 40325 23103
rect 40184 23072 40325 23100
rect 40184 23060 40190 23072
rect 40313 23069 40325 23072
rect 40359 23069 40371 23103
rect 40770 23100 40776 23112
rect 40731 23072 40776 23100
rect 40313 23063 40371 23069
rect 40770 23060 40776 23072
rect 40828 23060 40834 23112
rect 41046 23100 41052 23112
rect 41007 23072 41052 23100
rect 41046 23060 41052 23072
rect 41104 23060 41110 23112
rect 41598 23100 41604 23112
rect 41559 23072 41604 23100
rect 41598 23060 41604 23072
rect 41656 23060 41662 23112
rect 43806 23100 43812 23112
rect 43767 23072 43812 23100
rect 43806 23060 43812 23072
rect 43864 23060 43870 23112
rect 43898 23060 43904 23112
rect 43956 23100 43962 23112
rect 43993 23103 44051 23109
rect 43993 23100 44005 23103
rect 43956 23072 44005 23100
rect 43956 23060 43962 23072
rect 43993 23069 44005 23072
rect 44039 23069 44051 23103
rect 43993 23063 44051 23069
rect 44361 23103 44419 23109
rect 44361 23069 44373 23103
rect 44407 23069 44419 23103
rect 45646 23100 45652 23112
rect 45607 23072 45652 23100
rect 44361 23063 44419 23069
rect 40037 23035 40095 23041
rect 40037 23032 40049 23035
rect 40000 23004 40049 23032
rect 40000 22992 40006 23004
rect 40037 23001 40049 23004
rect 40083 23001 40095 23035
rect 40218 23032 40224 23044
rect 40179 23004 40224 23032
rect 40037 22995 40095 23001
rect 40218 22992 40224 23004
rect 40276 22992 40282 23044
rect 41064 23032 41092 23060
rect 41230 23032 41236 23044
rect 41064 23004 41236 23032
rect 41230 22992 41236 23004
rect 41288 23032 41294 23044
rect 44266 23032 44272 23044
rect 41288 23004 44272 23032
rect 41288 22992 41294 23004
rect 44266 22992 44272 23004
rect 44324 22992 44330 23044
rect 30607 22936 31064 22964
rect 30607 22933 30619 22936
rect 30561 22927 30619 22933
rect 31110 22924 31116 22976
rect 31168 22964 31174 22976
rect 32677 22967 32735 22973
rect 32677 22964 32689 22967
rect 31168 22936 32689 22964
rect 31168 22924 31174 22936
rect 32677 22933 32689 22936
rect 32723 22933 32735 22967
rect 37366 22964 37372 22976
rect 37327 22936 37372 22964
rect 32677 22927 32735 22933
rect 37366 22924 37372 22936
rect 37424 22924 37430 22976
rect 37458 22924 37464 22976
rect 37516 22964 37522 22976
rect 37737 22967 37795 22973
rect 37737 22964 37749 22967
rect 37516 22936 37749 22964
rect 37516 22924 37522 22936
rect 37737 22933 37749 22936
rect 37783 22933 37795 22967
rect 38378 22964 38384 22976
rect 38339 22936 38384 22964
rect 37737 22927 37795 22933
rect 38378 22924 38384 22936
rect 38436 22924 38442 22976
rect 40770 22964 40776 22976
rect 40731 22936 40776 22964
rect 40770 22924 40776 22936
rect 40828 22924 40834 22976
rect 44082 22924 44088 22976
rect 44140 22964 44146 22976
rect 44376 22964 44404 23063
rect 45646 23060 45652 23072
rect 45704 23060 45710 23112
rect 46474 23100 46480 23112
rect 46435 23072 46480 23100
rect 46474 23060 46480 23072
rect 46532 23060 46538 23112
rect 46661 23035 46719 23041
rect 46661 23001 46673 23035
rect 46707 23032 46719 23035
rect 47118 23032 47124 23044
rect 46707 23004 47124 23032
rect 46707 23001 46719 23004
rect 46661 22995 46719 23001
rect 47118 22992 47124 23004
rect 47176 22992 47182 23044
rect 48314 23032 48320 23044
rect 48275 23004 48320 23032
rect 48314 22992 48320 23004
rect 48372 22992 48378 23044
rect 44140 22936 44404 22964
rect 44140 22924 44146 22936
rect 44450 22924 44456 22976
rect 44508 22964 44514 22976
rect 44545 22967 44603 22973
rect 44545 22964 44557 22967
rect 44508 22936 44557 22964
rect 44508 22924 44514 22936
rect 44545 22933 44557 22936
rect 44591 22933 44603 22967
rect 44545 22927 44603 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 27062 22720 27068 22772
rect 27120 22760 27126 22772
rect 27341 22763 27399 22769
rect 27341 22760 27353 22763
rect 27120 22732 27353 22760
rect 27120 22720 27126 22732
rect 27341 22729 27353 22732
rect 27387 22729 27399 22763
rect 27614 22760 27620 22772
rect 27341 22723 27399 22729
rect 27540 22732 27620 22760
rect 2406 22652 2412 22704
rect 2464 22692 2470 22704
rect 5442 22692 5448 22704
rect 2464 22664 5448 22692
rect 2464 22652 2470 22664
rect 5442 22652 5448 22664
rect 5500 22692 5506 22704
rect 5500 22664 22094 22692
rect 5500 22652 5506 22664
rect 22066 22556 22094 22664
rect 23198 22624 23204 22636
rect 23159 22596 23204 22624
rect 23198 22584 23204 22596
rect 23256 22584 23262 22636
rect 23290 22584 23296 22636
rect 23348 22624 23354 22636
rect 23385 22627 23443 22633
rect 23385 22624 23397 22627
rect 23348 22596 23397 22624
rect 23348 22584 23354 22596
rect 23385 22593 23397 22596
rect 23431 22593 23443 22627
rect 26418 22624 26424 22636
rect 26379 22596 26424 22624
rect 23385 22587 23443 22593
rect 26418 22584 26424 22596
rect 26476 22584 26482 22636
rect 27540 22633 27568 22732
rect 27614 22720 27620 22732
rect 27672 22720 27678 22772
rect 28442 22760 28448 22772
rect 28403 22732 28448 22760
rect 28442 22720 28448 22732
rect 28500 22720 28506 22772
rect 36173 22763 36231 22769
rect 29748 22732 31754 22760
rect 29748 22692 29776 22732
rect 30466 22692 30472 22704
rect 28368 22664 29776 22692
rect 29840 22664 30472 22692
rect 27525 22627 27583 22633
rect 27525 22593 27537 22627
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 27614 22584 27620 22636
rect 27672 22624 27678 22636
rect 27893 22627 27951 22633
rect 27672 22596 27717 22624
rect 27672 22584 27678 22596
rect 27893 22593 27905 22627
rect 27939 22624 27951 22627
rect 28166 22624 28172 22636
rect 27939 22596 28172 22624
rect 27939 22593 27951 22596
rect 27893 22587 27951 22593
rect 28166 22584 28172 22596
rect 28224 22584 28230 22636
rect 28368 22633 28396 22664
rect 29840 22633 29868 22664
rect 30466 22652 30472 22664
rect 30524 22692 30530 22704
rect 30524 22664 30696 22692
rect 30524 22652 30530 22664
rect 28353 22627 28411 22633
rect 28353 22593 28365 22627
rect 28399 22593 28411 22627
rect 28353 22587 28411 22593
rect 29641 22627 29699 22633
rect 29641 22593 29653 22627
rect 29687 22593 29699 22627
rect 29641 22587 29699 22593
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 30374 22624 30380 22636
rect 30335 22596 30380 22624
rect 29825 22587 29883 22593
rect 28368 22556 28396 22587
rect 22066 22528 28396 22556
rect 26513 22491 26571 22497
rect 26513 22457 26525 22491
rect 26559 22488 26571 22491
rect 27522 22488 27528 22500
rect 26559 22460 27528 22488
rect 26559 22457 26571 22460
rect 26513 22451 26571 22457
rect 27522 22448 27528 22460
rect 27580 22448 27586 22500
rect 27798 22488 27804 22500
rect 27759 22460 27804 22488
rect 27798 22448 27804 22460
rect 27856 22448 27862 22500
rect 29656 22488 29684 22587
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 30668 22633 30696 22664
rect 30742 22652 30748 22704
rect 30800 22692 30806 22704
rect 31726 22692 31754 22732
rect 36173 22729 36185 22763
rect 36219 22760 36231 22763
rect 37458 22760 37464 22772
rect 36219 22732 37464 22760
rect 36219 22729 36231 22732
rect 36173 22723 36231 22729
rect 37458 22720 37464 22732
rect 37516 22720 37522 22772
rect 37550 22720 37556 22772
rect 37608 22760 37614 22772
rect 38105 22763 38163 22769
rect 38105 22760 38117 22763
rect 37608 22732 38117 22760
rect 37608 22720 37614 22732
rect 38105 22729 38117 22732
rect 38151 22729 38163 22763
rect 39669 22763 39727 22769
rect 38105 22723 38163 22729
rect 38626 22732 38980 22760
rect 36630 22692 36636 22704
rect 30800 22664 31524 22692
rect 31726 22664 36636 22692
rect 30800 22652 30806 22664
rect 31496 22636 31524 22664
rect 36630 22652 36636 22664
rect 36688 22652 36694 22704
rect 37366 22652 37372 22704
rect 37424 22692 37430 22704
rect 38626 22692 38654 22732
rect 37424 22664 38654 22692
rect 37424 22652 37430 22664
rect 30561 22627 30619 22633
rect 30561 22593 30573 22627
rect 30607 22593 30619 22627
rect 30561 22587 30619 22593
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22593 30711 22627
rect 30653 22587 30711 22593
rect 29914 22556 29920 22568
rect 29827 22528 29920 22556
rect 29914 22516 29920 22528
rect 29972 22556 29978 22568
rect 30576 22556 30604 22587
rect 30926 22584 30932 22636
rect 30984 22624 30990 22636
rect 31205 22627 31263 22633
rect 31205 22624 31217 22627
rect 30984 22596 31217 22624
rect 30984 22584 30990 22596
rect 31205 22593 31217 22596
rect 31251 22593 31263 22627
rect 31386 22624 31392 22636
rect 31347 22596 31392 22624
rect 31205 22587 31263 22593
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 31478 22584 31484 22636
rect 31536 22624 31542 22636
rect 31536 22596 31629 22624
rect 31536 22584 31542 22596
rect 33134 22584 33140 22636
rect 33192 22624 33198 22636
rect 33870 22633 33876 22636
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 33192 22596 33609 22624
rect 33192 22584 33198 22596
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 33864 22587 33876 22633
rect 33928 22624 33934 22636
rect 36354 22624 36360 22636
rect 33928 22596 33964 22624
rect 34992 22596 36360 22624
rect 33870 22584 33876 22587
rect 33928 22584 33934 22596
rect 31110 22556 31116 22568
rect 29972 22528 31116 22556
rect 29972 22516 29978 22528
rect 31110 22516 31116 22528
rect 31168 22516 31174 22568
rect 30377 22491 30435 22497
rect 30377 22488 30389 22491
rect 29656 22460 30389 22488
rect 30377 22457 30389 22460
rect 30423 22457 30435 22491
rect 30377 22451 30435 22457
rect 30650 22448 30656 22500
rect 30708 22488 30714 22500
rect 31205 22491 31263 22497
rect 31205 22488 31217 22491
rect 30708 22460 31217 22488
rect 30708 22448 30714 22460
rect 31205 22457 31217 22460
rect 31251 22457 31263 22491
rect 31205 22451 31263 22457
rect 23201 22423 23259 22429
rect 23201 22389 23213 22423
rect 23247 22420 23259 22423
rect 23382 22420 23388 22432
rect 23247 22392 23388 22420
rect 23247 22389 23259 22392
rect 23201 22383 23259 22389
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 29454 22420 29460 22432
rect 29415 22392 29460 22420
rect 29454 22380 29460 22392
rect 29512 22380 29518 22432
rect 30466 22380 30472 22432
rect 30524 22420 30530 22432
rect 32490 22420 32496 22432
rect 30524 22392 32496 22420
rect 30524 22380 30530 22392
rect 32490 22380 32496 22392
rect 32548 22380 32554 22432
rect 34698 22380 34704 22432
rect 34756 22420 34762 22432
rect 34992 22429 35020 22596
rect 36354 22584 36360 22596
rect 36412 22584 36418 22636
rect 36449 22627 36507 22633
rect 36449 22593 36461 22627
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 36262 22516 36268 22568
rect 36320 22556 36326 22568
rect 36464 22556 36492 22587
rect 36538 22584 36544 22636
rect 36596 22624 36602 22636
rect 36725 22627 36783 22633
rect 36725 22624 36737 22627
rect 36596 22596 36737 22624
rect 36596 22584 36602 22596
rect 36725 22593 36737 22596
rect 36771 22624 36783 22627
rect 37553 22627 37611 22633
rect 37553 22624 37565 22627
rect 36771 22596 37565 22624
rect 36771 22593 36783 22596
rect 36725 22587 36783 22593
rect 37553 22593 37565 22596
rect 37599 22593 37611 22627
rect 37734 22624 37740 22636
rect 37695 22596 37740 22624
rect 37553 22587 37611 22593
rect 37734 22584 37740 22596
rect 37792 22584 37798 22636
rect 37829 22627 37887 22633
rect 37829 22593 37841 22627
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 37921 22627 37979 22633
rect 37921 22593 37933 22627
rect 37967 22624 37979 22627
rect 38838 22624 38844 22636
rect 37967 22596 38844 22624
rect 37967 22593 37979 22596
rect 37921 22587 37979 22593
rect 36814 22556 36820 22568
rect 36320 22528 36820 22556
rect 36320 22516 36326 22528
rect 36814 22516 36820 22528
rect 36872 22516 36878 22568
rect 37844 22556 37872 22587
rect 38838 22584 38844 22596
rect 38896 22584 38902 22636
rect 38952 22633 38980 22732
rect 39669 22729 39681 22763
rect 39715 22760 39727 22763
rect 40034 22760 40040 22772
rect 39715 22732 40040 22760
rect 39715 22729 39727 22732
rect 39669 22723 39727 22729
rect 40034 22720 40040 22732
rect 40092 22720 40098 22772
rect 41509 22763 41567 22769
rect 41509 22729 41521 22763
rect 41555 22760 41567 22763
rect 41690 22760 41696 22772
rect 41555 22732 41696 22760
rect 41555 22729 41567 22732
rect 41509 22723 41567 22729
rect 41690 22720 41696 22732
rect 41748 22720 41754 22772
rect 43441 22763 43499 22769
rect 43441 22729 43453 22763
rect 43487 22760 43499 22763
rect 44082 22760 44088 22772
rect 43487 22732 44088 22760
rect 43487 22729 43499 22732
rect 43441 22723 43499 22729
rect 44082 22720 44088 22732
rect 44140 22760 44146 22772
rect 44269 22763 44327 22769
rect 44269 22760 44281 22763
rect 44140 22732 44281 22760
rect 44140 22720 44146 22732
rect 44269 22729 44281 22732
rect 44315 22729 44327 22763
rect 47118 22760 47124 22772
rect 47079 22732 47124 22760
rect 44269 22723 44327 22729
rect 47118 22720 47124 22732
rect 47176 22720 47182 22772
rect 41598 22692 41604 22704
rect 40144 22664 41604 22692
rect 38933 22627 38991 22633
rect 38933 22593 38945 22627
rect 38979 22593 38991 22627
rect 39114 22624 39120 22636
rect 39075 22596 39120 22624
rect 38933 22587 38991 22593
rect 39114 22584 39120 22596
rect 39172 22584 39178 22636
rect 39298 22624 39304 22636
rect 39259 22596 39304 22624
rect 39298 22584 39304 22596
rect 39356 22584 39362 22636
rect 39482 22624 39488 22636
rect 39443 22596 39488 22624
rect 39482 22584 39488 22596
rect 39540 22584 39546 22636
rect 40144 22633 40172 22664
rect 41598 22652 41604 22664
rect 41656 22652 41662 22704
rect 44174 22692 44180 22704
rect 44135 22664 44180 22692
rect 44174 22652 44180 22664
rect 44232 22652 44238 22704
rect 44637 22695 44695 22701
rect 44637 22661 44649 22695
rect 44683 22692 44695 22695
rect 45370 22692 45376 22704
rect 44683 22664 45376 22692
rect 44683 22661 44695 22664
rect 44637 22655 44695 22661
rect 45370 22652 45376 22664
rect 45428 22652 45434 22704
rect 46474 22652 46480 22704
rect 46532 22692 46538 22704
rect 46532 22664 47992 22692
rect 46532 22652 46538 22664
rect 40129 22627 40187 22633
rect 40129 22593 40141 22627
rect 40175 22593 40187 22627
rect 40129 22587 40187 22593
rect 40396 22627 40454 22633
rect 40396 22593 40408 22627
rect 40442 22624 40454 22627
rect 40770 22624 40776 22636
rect 40442 22596 40776 22624
rect 40442 22593 40454 22596
rect 40396 22587 40454 22593
rect 40770 22584 40776 22596
rect 40828 22584 40834 22636
rect 43346 22624 43352 22636
rect 43307 22596 43352 22624
rect 43346 22584 43352 22596
rect 43404 22584 43410 22636
rect 44450 22624 44456 22636
rect 44411 22596 44456 22624
rect 44450 22584 44456 22596
rect 44508 22584 44514 22636
rect 45094 22624 45100 22636
rect 45055 22596 45100 22624
rect 45094 22584 45100 22596
rect 45152 22584 45158 22636
rect 47026 22624 47032 22636
rect 46987 22596 47032 22624
rect 47026 22584 47032 22596
rect 47084 22584 47090 22636
rect 47964 22633 47992 22664
rect 47949 22627 48007 22633
rect 47949 22593 47961 22627
rect 47995 22593 48007 22627
rect 47949 22587 48007 22593
rect 39022 22556 39028 22568
rect 37844 22528 39028 22556
rect 39022 22516 39028 22528
rect 39080 22556 39086 22568
rect 39209 22559 39267 22565
rect 39209 22556 39221 22559
rect 39080 22528 39221 22556
rect 39080 22516 39086 22528
rect 39209 22525 39221 22528
rect 39255 22525 39267 22559
rect 39209 22519 39267 22525
rect 44266 22516 44272 22568
rect 44324 22556 44330 22568
rect 44545 22559 44603 22565
rect 44545 22556 44557 22559
rect 44324 22528 44557 22556
rect 44324 22516 44330 22528
rect 44545 22525 44557 22528
rect 44591 22525 44603 22559
rect 44545 22519 44603 22525
rect 36633 22491 36691 22497
rect 36633 22457 36645 22491
rect 36679 22488 36691 22491
rect 37734 22488 37740 22500
rect 36679 22460 37740 22488
rect 36679 22457 36691 22460
rect 36633 22451 36691 22457
rect 37734 22448 37740 22460
rect 37792 22448 37798 22500
rect 43990 22448 43996 22500
rect 44048 22488 44054 22500
rect 45189 22491 45247 22497
rect 45189 22488 45201 22491
rect 44048 22460 45201 22488
rect 44048 22448 44054 22460
rect 45189 22457 45201 22460
rect 45235 22457 45247 22491
rect 45189 22451 45247 22457
rect 34977 22423 35035 22429
rect 34977 22420 34989 22423
rect 34756 22392 34989 22420
rect 34756 22380 34762 22392
rect 34977 22389 34989 22392
rect 35023 22389 35035 22423
rect 34977 22383 35035 22389
rect 41506 22380 41512 22432
rect 41564 22420 41570 22432
rect 45646 22420 45652 22432
rect 41564 22392 45652 22420
rect 41564 22380 41570 22392
rect 45646 22380 45652 22392
rect 45704 22380 45710 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 26970 22176 26976 22228
rect 27028 22216 27034 22228
rect 30374 22216 30380 22228
rect 27028 22188 30380 22216
rect 27028 22176 27034 22188
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 31110 22216 31116 22228
rect 31071 22188 31116 22216
rect 31110 22176 31116 22188
rect 31168 22176 31174 22228
rect 33870 22176 33876 22228
rect 33928 22216 33934 22228
rect 34057 22219 34115 22225
rect 34057 22216 34069 22219
rect 33928 22188 34069 22216
rect 33928 22176 33934 22188
rect 34057 22185 34069 22188
rect 34103 22185 34115 22219
rect 34057 22179 34115 22185
rect 36630 22176 36636 22228
rect 36688 22216 36694 22228
rect 41506 22216 41512 22228
rect 36688 22188 41512 22216
rect 36688 22176 36694 22188
rect 41506 22176 41512 22188
rect 41564 22176 41570 22228
rect 41598 22176 41604 22228
rect 41656 22216 41662 22228
rect 42702 22216 42708 22228
rect 41656 22188 42708 22216
rect 41656 22176 41662 22188
rect 42702 22176 42708 22188
rect 42760 22176 42766 22228
rect 42981 22219 43039 22225
rect 42981 22185 42993 22219
rect 43027 22216 43039 22219
rect 43346 22216 43352 22228
rect 43027 22188 43352 22216
rect 43027 22185 43039 22188
rect 42981 22179 43039 22185
rect 34149 22151 34207 22157
rect 34149 22117 34161 22151
rect 34195 22148 34207 22151
rect 34885 22151 34943 22157
rect 34885 22148 34897 22151
rect 34195 22120 34897 22148
rect 34195 22117 34207 22120
rect 34149 22111 34207 22117
rect 34885 22117 34897 22120
rect 34931 22117 34943 22151
rect 34885 22111 34943 22117
rect 2774 22080 2780 22092
rect 2735 22052 2780 22080
rect 2774 22040 2780 22052
rect 2832 22040 2838 22092
rect 23109 22083 23167 22089
rect 23109 22049 23121 22083
rect 23155 22080 23167 22083
rect 26234 22080 26240 22092
rect 23155 22052 26240 22080
rect 23155 22049 23167 22052
rect 23109 22043 23167 22049
rect 26234 22040 26240 22052
rect 26292 22040 26298 22092
rect 34790 22080 34796 22092
rect 34072 22052 34796 22080
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 22830 21972 22836 22024
rect 22888 22012 22894 22024
rect 23198 22012 23204 22024
rect 22888 21984 23204 22012
rect 22888 21972 22894 21984
rect 23198 21972 23204 21984
rect 23256 22012 23262 22024
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 23256 21984 23305 22012
rect 23256 21972 23262 21984
rect 23293 21981 23305 21984
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 21981 23627 22015
rect 29730 22012 29736 22024
rect 29691 21984 29736 22012
rect 23569 21975 23627 21981
rect 1762 21944 1768 21956
rect 1723 21916 1768 21944
rect 1762 21904 1768 21916
rect 1820 21904 1826 21956
rect 23584 21944 23612 21975
rect 29730 21972 29736 21984
rect 29788 21972 29794 22024
rect 34072 22021 34100 22052
rect 34790 22040 34796 22052
rect 34848 22040 34854 22092
rect 34057 22015 34115 22021
rect 34057 21981 34069 22015
rect 34103 21981 34115 22015
rect 34057 21975 34115 21981
rect 34698 21972 34704 22024
rect 34756 22012 34762 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34756 21984 34897 22012
rect 34756 21972 34762 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 35161 22015 35219 22021
rect 35161 21981 35173 22015
rect 35207 22012 35219 22015
rect 35342 22012 35348 22024
rect 35207 21984 35348 22012
rect 35207 21981 35219 21984
rect 35161 21975 35219 21981
rect 35342 21972 35348 21984
rect 35400 21972 35406 22024
rect 37274 22012 37280 22024
rect 37235 21984 37280 22012
rect 37274 21972 37280 21984
rect 37332 21972 37338 22024
rect 40494 21972 40500 22024
rect 40552 22012 40558 22024
rect 40957 22015 41015 22021
rect 40957 22012 40969 22015
rect 40552 21984 40969 22012
rect 40552 21972 40558 21984
rect 40957 21981 40969 21984
rect 41003 21981 41015 22015
rect 40957 21975 41015 21981
rect 41138 21972 41144 22024
rect 41196 22012 41202 22024
rect 41598 22012 41604 22024
rect 41196 21984 41414 22012
rect 41559 21984 41604 22012
rect 41196 21972 41202 21984
rect 23216 21916 23612 21944
rect 23216 21888 23244 21916
rect 29454 21904 29460 21956
rect 29512 21944 29518 21956
rect 29978 21947 30036 21953
rect 29978 21944 29990 21947
rect 29512 21916 29990 21944
rect 29512 21904 29518 21916
rect 29978 21913 29990 21916
rect 30024 21913 30036 21947
rect 29978 21907 30036 21913
rect 33962 21904 33968 21956
rect 34020 21944 34026 21956
rect 34330 21944 34336 21956
rect 34020 21916 34336 21944
rect 34020 21904 34026 21916
rect 34330 21904 34336 21916
rect 34388 21904 34394 21956
rect 34606 21904 34612 21956
rect 34664 21944 34670 21956
rect 35069 21947 35127 21953
rect 35069 21944 35081 21947
rect 34664 21916 35081 21944
rect 34664 21904 34670 21916
rect 35069 21913 35081 21916
rect 35115 21913 35127 21947
rect 35069 21907 35127 21913
rect 37544 21947 37602 21953
rect 37544 21913 37556 21947
rect 37590 21944 37602 21947
rect 38378 21944 38384 21956
rect 37590 21916 38384 21944
rect 37590 21913 37602 21916
rect 37544 21907 37602 21913
rect 38378 21904 38384 21916
rect 38436 21904 38442 21956
rect 41386 21944 41414 21984
rect 41598 21972 41604 21984
rect 41656 21972 41662 22024
rect 42996 22012 43024 22179
rect 43346 22176 43352 22188
rect 43404 22176 43410 22228
rect 43990 22080 43996 22092
rect 43951 22052 43996 22080
rect 43990 22040 43996 22052
rect 44048 22040 44054 22092
rect 41708 21984 43024 22012
rect 43901 22015 43959 22021
rect 41708 21944 41736 21984
rect 43901 21981 43913 22015
rect 43947 22012 43959 22015
rect 44082 22012 44088 22024
rect 43947 21984 44088 22012
rect 43947 21981 43959 21984
rect 43901 21975 43959 21981
rect 44082 21972 44088 21984
rect 44140 21972 44146 22024
rect 46474 22012 46480 22024
rect 46435 21984 46480 22012
rect 46474 21972 46480 21984
rect 46532 21972 46538 22024
rect 41386 21916 41736 21944
rect 41868 21947 41926 21953
rect 41868 21913 41880 21947
rect 41914 21944 41926 21947
rect 42058 21944 42064 21956
rect 41914 21916 42064 21944
rect 41914 21913 41926 21916
rect 41868 21907 41926 21913
rect 42058 21904 42064 21916
rect 42116 21904 42122 21956
rect 46661 21947 46719 21953
rect 46661 21913 46673 21947
rect 46707 21944 46719 21947
rect 47118 21944 47124 21956
rect 46707 21916 47124 21944
rect 46707 21913 46719 21916
rect 46661 21907 46719 21913
rect 47118 21904 47124 21916
rect 47176 21904 47182 21956
rect 48314 21944 48320 21956
rect 48275 21916 48320 21944
rect 48314 21904 48320 21916
rect 48372 21904 48378 21956
rect 23198 21836 23204 21888
rect 23256 21836 23262 21888
rect 23382 21836 23388 21888
rect 23440 21876 23446 21888
rect 23477 21879 23535 21885
rect 23477 21876 23489 21879
rect 23440 21848 23489 21876
rect 23440 21836 23446 21848
rect 23477 21845 23489 21848
rect 23523 21845 23535 21879
rect 23477 21839 23535 21845
rect 37734 21836 37740 21888
rect 37792 21876 37798 21888
rect 38657 21879 38715 21885
rect 38657 21876 38669 21879
rect 37792 21848 38669 21876
rect 37792 21836 37798 21848
rect 38657 21845 38669 21848
rect 38703 21845 38715 21879
rect 38657 21839 38715 21845
rect 41049 21879 41107 21885
rect 41049 21845 41061 21879
rect 41095 21876 41107 21879
rect 41782 21876 41788 21888
rect 41095 21848 41788 21876
rect 41095 21845 41107 21848
rect 41049 21839 41107 21845
rect 41782 21836 41788 21848
rect 41840 21836 41846 21888
rect 44174 21836 44180 21888
rect 44232 21876 44238 21888
rect 44269 21879 44327 21885
rect 44269 21876 44281 21879
rect 44232 21848 44281 21876
rect 44232 21836 44238 21848
rect 44269 21845 44281 21848
rect 44315 21845 44327 21879
rect 44269 21839 44327 21845
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1762 21632 1768 21684
rect 1820 21672 1826 21684
rect 2869 21675 2927 21681
rect 2869 21672 2881 21675
rect 1820 21644 2881 21672
rect 1820 21632 1826 21644
rect 2869 21641 2881 21644
rect 2915 21641 2927 21675
rect 22830 21672 22836 21684
rect 22791 21644 22836 21672
rect 2869 21635 2927 21641
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 23474 21672 23480 21684
rect 22940 21644 23480 21672
rect 22940 21604 22968 21644
rect 23474 21632 23480 21644
rect 23532 21672 23538 21684
rect 25777 21675 25835 21681
rect 25777 21672 25789 21675
rect 23532 21644 25789 21672
rect 23532 21632 23538 21644
rect 25777 21641 25789 21644
rect 25823 21672 25835 21675
rect 26418 21672 26424 21684
rect 25823 21644 26424 21672
rect 25823 21641 25835 21644
rect 25777 21635 25835 21641
rect 26418 21632 26424 21644
rect 26476 21632 26482 21684
rect 30009 21675 30067 21681
rect 30009 21641 30021 21675
rect 30055 21672 30067 21675
rect 30190 21672 30196 21684
rect 30055 21644 30196 21672
rect 30055 21641 30067 21644
rect 30009 21635 30067 21641
rect 30190 21632 30196 21644
rect 30248 21672 30254 21684
rect 31386 21672 31392 21684
rect 30248 21644 31392 21672
rect 30248 21632 30254 21644
rect 31386 21632 31392 21644
rect 31444 21632 31450 21684
rect 37829 21675 37887 21681
rect 37829 21641 37841 21675
rect 37875 21672 37887 21675
rect 38470 21672 38476 21684
rect 37875 21644 38476 21672
rect 37875 21641 37887 21644
rect 37829 21635 37887 21641
rect 38470 21632 38476 21644
rect 38528 21632 38534 21684
rect 44453 21675 44511 21681
rect 44453 21672 44465 21675
rect 41616 21644 44465 21672
rect 22572 21576 22968 21604
rect 29825 21607 29883 21613
rect 1578 21496 1584 21548
rect 1636 21536 1642 21548
rect 2317 21539 2375 21545
rect 2317 21536 2329 21539
rect 1636 21508 2329 21536
rect 1636 21496 1642 21508
rect 2317 21505 2329 21508
rect 2363 21505 2375 21539
rect 2317 21499 2375 21505
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21536 2835 21539
rect 2958 21536 2964 21548
rect 2823 21508 2964 21536
rect 2823 21505 2835 21508
rect 2777 21499 2835 21505
rect 2958 21496 2964 21508
rect 3016 21496 3022 21548
rect 22572 21545 22600 21576
rect 29825 21573 29837 21607
rect 29871 21604 29883 21607
rect 30466 21604 30472 21616
rect 29871 21576 30472 21604
rect 29871 21573 29883 21576
rect 29825 21567 29883 21573
rect 30466 21564 30472 21576
rect 30524 21564 30530 21616
rect 41616 21613 41644 21644
rect 44453 21641 44465 21644
rect 44499 21641 44511 21675
rect 47118 21672 47124 21684
rect 47079 21644 47124 21672
rect 44453 21635 44511 21641
rect 47118 21632 47124 21644
rect 47176 21632 47182 21684
rect 41601 21607 41659 21613
rect 41601 21573 41613 21607
rect 41647 21573 41659 21607
rect 42058 21604 42064 21616
rect 42019 21576 42064 21604
rect 41601 21567 41659 21573
rect 42058 21564 42064 21576
rect 42116 21564 42122 21616
rect 46474 21564 46480 21616
rect 46532 21604 46538 21616
rect 46532 21576 47992 21604
rect 46532 21564 46538 21576
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21536 22707 21539
rect 23106 21536 23112 21548
rect 22695 21508 23112 21536
rect 22695 21505 22707 21508
rect 22649 21499 22707 21505
rect 23106 21496 23112 21508
rect 23164 21496 23170 21548
rect 23474 21496 23480 21548
rect 23532 21545 23538 21548
rect 23532 21539 23581 21545
rect 23532 21505 23535 21539
rect 23569 21505 23581 21539
rect 23532 21499 23581 21505
rect 23658 21542 23716 21548
rect 23658 21508 23670 21542
rect 23704 21508 23716 21542
rect 23658 21502 23716 21508
rect 23532 21496 23538 21499
rect 23676 21468 23704 21502
rect 23750 21496 23756 21548
rect 23808 21536 23814 21548
rect 23937 21539 23995 21545
rect 23808 21508 23853 21536
rect 23808 21496 23814 21508
rect 23937 21505 23949 21539
rect 23983 21536 23995 21539
rect 24026 21536 24032 21548
rect 23983 21508 24032 21536
rect 23983 21505 23995 21508
rect 23937 21499 23995 21505
rect 24026 21496 24032 21508
rect 24084 21496 24090 21548
rect 24394 21536 24400 21548
rect 24355 21508 24400 21536
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 24653 21539 24711 21545
rect 24653 21536 24665 21539
rect 24504 21508 24665 21536
rect 24504 21468 24532 21508
rect 24653 21505 24665 21508
rect 24699 21505 24711 21539
rect 24653 21499 24711 21505
rect 26878 21496 26884 21548
rect 26936 21536 26942 21548
rect 27525 21539 27583 21545
rect 27525 21536 27537 21539
rect 26936 21508 27537 21536
rect 26936 21496 26942 21508
rect 27525 21505 27537 21508
rect 27571 21505 27583 21539
rect 27525 21499 27583 21505
rect 27709 21539 27767 21545
rect 27709 21505 27721 21539
rect 27755 21536 27767 21539
rect 28258 21536 28264 21548
rect 27755 21508 28264 21536
rect 27755 21505 27767 21508
rect 27709 21499 27767 21505
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 30101 21539 30159 21545
rect 30101 21505 30113 21539
rect 30147 21536 30159 21539
rect 31478 21536 31484 21548
rect 30147 21508 31484 21536
rect 30147 21505 30159 21508
rect 30101 21499 30159 21505
rect 31478 21496 31484 21508
rect 31536 21496 31542 21548
rect 37642 21536 37648 21548
rect 37603 21508 37648 21536
rect 37642 21496 37648 21508
rect 37700 21496 37706 21548
rect 41690 21536 41696 21548
rect 41651 21508 41696 21536
rect 41690 21496 41696 21508
rect 41748 21496 41754 21548
rect 41782 21496 41788 21548
rect 41840 21536 41846 21548
rect 41877 21539 41935 21545
rect 41877 21536 41889 21539
rect 41840 21508 41889 21536
rect 41840 21496 41846 21508
rect 41877 21505 41889 21508
rect 41923 21505 41935 21539
rect 41877 21499 41935 21505
rect 44085 21539 44143 21545
rect 44085 21505 44097 21539
rect 44131 21536 44143 21539
rect 44266 21536 44272 21548
rect 44131 21508 44272 21536
rect 44131 21505 44143 21508
rect 44085 21499 44143 21505
rect 44266 21496 44272 21508
rect 44324 21496 44330 21548
rect 47026 21536 47032 21548
rect 46987 21508 47032 21536
rect 47026 21496 47032 21508
rect 47084 21496 47090 21548
rect 47964 21545 47992 21576
rect 47949 21539 48007 21545
rect 47949 21505 47961 21539
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 23676 21440 23796 21468
rect 2314 21360 2320 21412
rect 2372 21400 2378 21412
rect 2682 21400 2688 21412
rect 2372 21372 2688 21400
rect 2372 21360 2378 21372
rect 2682 21360 2688 21372
rect 2740 21360 2746 21412
rect 23293 21403 23351 21409
rect 23293 21369 23305 21403
rect 23339 21369 23351 21403
rect 23768 21400 23796 21440
rect 24412 21440 24532 21468
rect 37461 21471 37519 21477
rect 23842 21400 23848 21412
rect 23768 21372 23848 21400
rect 23293 21363 23351 21369
rect 23308 21332 23336 21363
rect 23842 21360 23848 21372
rect 23900 21360 23906 21412
rect 24412 21332 24440 21440
rect 37461 21437 37473 21471
rect 37507 21468 37519 21471
rect 37734 21468 37740 21480
rect 37507 21440 37740 21468
rect 37507 21437 37519 21440
rect 37461 21431 37519 21437
rect 37734 21428 37740 21440
rect 37792 21428 37798 21480
rect 41414 21428 41420 21480
rect 41472 21468 41478 21480
rect 41969 21471 42027 21477
rect 41969 21468 41981 21471
rect 41472 21440 41981 21468
rect 41472 21428 41478 21440
rect 41969 21437 41981 21440
rect 42015 21437 42027 21471
rect 44174 21468 44180 21480
rect 44135 21440 44180 21468
rect 41969 21431 42027 21437
rect 44174 21428 44180 21440
rect 44232 21428 44238 21480
rect 23308 21304 24440 21332
rect 27430 21292 27436 21344
rect 27488 21332 27494 21344
rect 27525 21335 27583 21341
rect 27525 21332 27537 21335
rect 27488 21304 27537 21332
rect 27488 21292 27494 21304
rect 27525 21301 27537 21304
rect 27571 21301 27583 21335
rect 27525 21295 27583 21301
rect 29825 21335 29883 21341
rect 29825 21301 29837 21335
rect 29871 21332 29883 21335
rect 29914 21332 29920 21344
rect 29871 21304 29920 21332
rect 29871 21301 29883 21304
rect 29825 21295 29883 21301
rect 29914 21292 29920 21304
rect 29972 21292 29978 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 23750 21088 23756 21140
rect 23808 21128 23814 21140
rect 24673 21131 24731 21137
rect 24673 21128 24685 21131
rect 23808 21100 24685 21128
rect 23808 21088 23814 21100
rect 24673 21097 24685 21100
rect 24719 21097 24731 21131
rect 28258 21128 28264 21140
rect 28219 21100 28264 21128
rect 24673 21091 24731 21097
rect 28258 21088 28264 21100
rect 28316 21088 28322 21140
rect 31113 21131 31171 21137
rect 31113 21097 31125 21131
rect 31159 21128 31171 21131
rect 31386 21128 31392 21140
rect 31159 21100 31392 21128
rect 31159 21097 31171 21100
rect 31113 21091 31171 21097
rect 31386 21088 31392 21100
rect 31444 21088 31450 21140
rect 31478 21088 31484 21140
rect 31536 21128 31542 21140
rect 32953 21131 33011 21137
rect 32953 21128 32965 21131
rect 31536 21100 32965 21128
rect 31536 21088 31542 21100
rect 32953 21097 32965 21100
rect 32999 21097 33011 21131
rect 44634 21128 44640 21140
rect 44547 21100 44640 21128
rect 32953 21091 33011 21097
rect 44634 21088 44640 21100
rect 44692 21128 44698 21140
rect 45094 21128 45100 21140
rect 44692 21100 45100 21128
rect 44692 21088 44698 21100
rect 45094 21088 45100 21100
rect 45152 21088 45158 21140
rect 23106 21020 23112 21072
rect 23164 21060 23170 21072
rect 23164 21032 23336 21060
rect 23164 21020 23170 21032
rect 23198 20992 23204 21004
rect 23159 20964 23204 20992
rect 23198 20952 23204 20964
rect 23256 20952 23262 21004
rect 23308 20992 23336 21032
rect 24394 21020 24400 21072
rect 24452 21060 24458 21072
rect 24452 21032 26924 21060
rect 24452 21020 24458 21032
rect 26896 21001 26924 21032
rect 25961 20995 26019 21001
rect 25961 20992 25973 20995
rect 23308 20964 25973 20992
rect 25961 20961 25973 20964
rect 26007 20961 26019 20995
rect 25961 20955 26019 20961
rect 26881 20995 26939 21001
rect 26881 20961 26893 20995
rect 26927 20961 26939 20995
rect 26881 20955 26939 20961
rect 2038 20884 2044 20936
rect 2096 20924 2102 20936
rect 2317 20927 2375 20933
rect 2317 20924 2329 20927
rect 2096 20896 2329 20924
rect 2096 20884 2102 20896
rect 2317 20893 2329 20896
rect 2363 20893 2375 20927
rect 2317 20887 2375 20893
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 23382 20924 23388 20936
rect 23155 20896 23388 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 23382 20884 23388 20896
rect 23440 20884 23446 20936
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 23492 20896 24593 20924
rect 23492 20797 23520 20896
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 26053 20927 26111 20933
rect 26053 20893 26065 20927
rect 26099 20924 26111 20927
rect 26896 20924 26924 20955
rect 42702 20952 42708 21004
rect 42760 20992 42766 21004
rect 43257 20995 43315 21001
rect 43257 20992 43269 20995
rect 42760 20964 43269 20992
rect 42760 20952 42766 20964
rect 43257 20961 43269 20964
rect 43303 20961 43315 20995
rect 43257 20955 43315 20961
rect 29730 20924 29736 20936
rect 26099 20896 26832 20924
rect 26896 20896 29736 20924
rect 26099 20893 26111 20896
rect 26053 20887 26111 20893
rect 23842 20816 23848 20868
rect 23900 20856 23906 20868
rect 24780 20856 24808 20887
rect 25314 20856 25320 20868
rect 23900 20828 25320 20856
rect 23900 20816 23906 20828
rect 25314 20816 25320 20828
rect 25372 20856 25378 20868
rect 26694 20856 26700 20868
rect 25372 20828 26700 20856
rect 25372 20816 25378 20828
rect 26694 20816 26700 20828
rect 26752 20816 26758 20868
rect 23477 20791 23535 20797
rect 23477 20757 23489 20791
rect 23523 20757 23535 20791
rect 23477 20751 23535 20757
rect 26326 20748 26332 20800
rect 26384 20788 26390 20800
rect 26421 20791 26479 20797
rect 26421 20788 26433 20791
rect 26384 20760 26433 20788
rect 26384 20748 26390 20760
rect 26421 20757 26433 20760
rect 26467 20757 26479 20791
rect 26804 20788 26832 20896
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 31294 20884 31300 20936
rect 31352 20924 31358 20936
rect 31573 20927 31631 20933
rect 31573 20924 31585 20927
rect 31352 20896 31585 20924
rect 31352 20884 31358 20896
rect 31573 20893 31585 20896
rect 31619 20924 31631 20927
rect 32306 20924 32312 20936
rect 31619 20896 32312 20924
rect 31619 20893 31631 20896
rect 31573 20887 31631 20893
rect 32306 20884 32312 20896
rect 32364 20924 32370 20936
rect 33042 20924 33048 20936
rect 32364 20896 33048 20924
rect 32364 20884 32370 20896
rect 33042 20884 33048 20896
rect 33100 20924 33106 20936
rect 34885 20927 34943 20933
rect 34885 20924 34897 20927
rect 33100 20896 34897 20924
rect 33100 20884 33106 20896
rect 34885 20893 34897 20896
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 27148 20859 27206 20865
rect 27148 20825 27160 20859
rect 27194 20856 27206 20859
rect 27522 20856 27528 20868
rect 27194 20828 27528 20856
rect 27194 20825 27206 20828
rect 27148 20819 27206 20825
rect 27522 20816 27528 20828
rect 27580 20816 27586 20868
rect 29822 20816 29828 20868
rect 29880 20856 29886 20868
rect 31846 20865 31852 20868
rect 29978 20859 30036 20865
rect 29978 20856 29990 20859
rect 29880 20828 29990 20856
rect 29880 20816 29886 20828
rect 29978 20825 29990 20828
rect 30024 20825 30036 20859
rect 29978 20819 30036 20825
rect 31840 20819 31852 20865
rect 31904 20856 31910 20868
rect 35152 20859 35210 20865
rect 31904 20828 31940 20856
rect 31846 20816 31852 20819
rect 31904 20816 31910 20828
rect 35152 20825 35164 20859
rect 35198 20856 35210 20859
rect 35342 20856 35348 20868
rect 35198 20828 35348 20856
rect 35198 20825 35210 20828
rect 35152 20819 35210 20825
rect 35342 20816 35348 20828
rect 35400 20816 35406 20868
rect 42978 20816 42984 20868
rect 43036 20856 43042 20868
rect 43502 20859 43560 20865
rect 43502 20856 43514 20859
rect 43036 20828 43514 20856
rect 43036 20816 43042 20828
rect 43502 20825 43514 20828
rect 43548 20825 43560 20859
rect 43502 20819 43560 20825
rect 28166 20788 28172 20800
rect 26804 20760 28172 20788
rect 26421 20751 26479 20757
rect 28166 20748 28172 20760
rect 28224 20748 28230 20800
rect 36262 20788 36268 20800
rect 36223 20760 36268 20788
rect 36262 20748 36268 20760
rect 36320 20748 36326 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 23290 20584 23296 20596
rect 23251 20556 23296 20584
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 26605 20587 26663 20593
rect 26605 20553 26617 20587
rect 26651 20553 26663 20587
rect 26605 20547 26663 20553
rect 26620 20516 26648 20547
rect 26694 20544 26700 20596
rect 26752 20584 26758 20596
rect 27249 20587 27307 20593
rect 27249 20584 27261 20587
rect 26752 20556 27261 20584
rect 26752 20544 26758 20556
rect 27249 20553 27261 20556
rect 27295 20553 27307 20587
rect 28166 20584 28172 20596
rect 28127 20556 28172 20584
rect 27249 20547 27307 20553
rect 28166 20544 28172 20556
rect 28224 20544 28230 20596
rect 29733 20587 29791 20593
rect 29733 20553 29745 20587
rect 29779 20584 29791 20587
rect 29822 20584 29828 20596
rect 29779 20556 29828 20584
rect 29779 20553 29791 20556
rect 29733 20547 29791 20553
rect 29822 20544 29828 20556
rect 29880 20544 29886 20596
rect 31665 20587 31723 20593
rect 31665 20553 31677 20587
rect 31711 20584 31723 20587
rect 31846 20584 31852 20596
rect 31711 20556 31852 20584
rect 31711 20553 31723 20556
rect 31665 20547 31723 20553
rect 31846 20544 31852 20556
rect 31904 20544 31910 20596
rect 35342 20584 35348 20596
rect 35303 20556 35348 20584
rect 35342 20544 35348 20556
rect 35400 20544 35406 20596
rect 35636 20556 37964 20584
rect 27157 20519 27215 20525
rect 27157 20516 27169 20519
rect 26620 20488 27169 20516
rect 27157 20485 27169 20488
rect 27203 20485 27215 20519
rect 34330 20516 34336 20528
rect 27157 20479 27215 20485
rect 31772 20488 34336 20516
rect 2038 20448 2044 20460
rect 1999 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 23106 20408 23112 20460
rect 23164 20448 23170 20460
rect 23201 20451 23259 20457
rect 23201 20448 23213 20451
rect 23164 20420 23213 20448
rect 23164 20408 23170 20420
rect 23201 20417 23213 20420
rect 23247 20417 23259 20451
rect 23201 20411 23259 20417
rect 23385 20451 23443 20457
rect 23385 20417 23397 20451
rect 23431 20448 23443 20451
rect 23474 20448 23480 20460
rect 23431 20420 23480 20448
rect 23431 20417 23443 20420
rect 23385 20411 23443 20417
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 26234 20448 26240 20460
rect 26195 20420 26240 20448
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 27430 20448 27436 20460
rect 27391 20420 27436 20448
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 28077 20451 28135 20457
rect 28077 20417 28089 20451
rect 28123 20448 28135 20451
rect 28258 20448 28264 20460
rect 28123 20420 28264 20448
rect 28123 20417 28135 20420
rect 28077 20411 28135 20417
rect 28258 20408 28264 20420
rect 28316 20408 28322 20460
rect 29914 20448 29920 20460
rect 29875 20420 29920 20448
rect 29914 20408 29920 20420
rect 29972 20408 29978 20460
rect 30190 20448 30196 20460
rect 30151 20420 30196 20448
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 31478 20408 31484 20460
rect 31536 20448 31542 20460
rect 31772 20457 31800 20488
rect 34330 20476 34336 20488
rect 34388 20476 34394 20528
rect 35636 20516 35664 20556
rect 34440 20488 35664 20516
rect 37936 20516 37964 20556
rect 38470 20544 38476 20596
rect 38528 20584 38534 20596
rect 42978 20584 42984 20596
rect 38528 20556 42564 20584
rect 42939 20556 42984 20584
rect 38528 20544 38534 20556
rect 38194 20516 38200 20528
rect 37936 20488 38200 20516
rect 31573 20451 31631 20457
rect 31573 20448 31585 20451
rect 31536 20420 31585 20448
rect 31536 20408 31542 20420
rect 31573 20417 31585 20420
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20417 31815 20451
rect 32306 20448 32312 20460
rect 32267 20420 32312 20448
rect 31757 20411 31815 20417
rect 32306 20408 32312 20420
rect 32364 20408 32370 20460
rect 32576 20451 32634 20457
rect 32576 20417 32588 20451
rect 32622 20448 32634 20451
rect 32858 20448 32864 20460
rect 32622 20420 32864 20448
rect 32622 20417 32634 20420
rect 32576 20411 32634 20417
rect 32858 20408 32864 20420
rect 32916 20408 32922 20460
rect 33870 20408 33876 20460
rect 33928 20448 33934 20460
rect 34440 20448 34468 20488
rect 34606 20448 34612 20460
rect 33928 20420 34468 20448
rect 34567 20420 34612 20448
rect 33928 20408 33934 20420
rect 34606 20408 34612 20420
rect 34664 20408 34670 20460
rect 34790 20448 34796 20460
rect 34751 20420 34796 20448
rect 34790 20408 34796 20420
rect 34848 20408 34854 20460
rect 34992 20457 35020 20488
rect 38194 20476 38200 20488
rect 38252 20476 38258 20528
rect 41598 20516 41604 20528
rect 40512 20488 41604 20516
rect 34977 20451 35035 20457
rect 34977 20417 34989 20451
rect 35023 20417 35035 20451
rect 34977 20411 35035 20417
rect 35161 20451 35219 20457
rect 35161 20417 35173 20451
rect 35207 20417 35219 20451
rect 35802 20448 35808 20460
rect 35763 20420 35808 20448
rect 35161 20411 35219 20417
rect 2225 20383 2283 20389
rect 2225 20349 2237 20383
rect 2271 20380 2283 20383
rect 2498 20380 2504 20392
rect 2271 20352 2504 20380
rect 2271 20349 2283 20352
rect 2225 20343 2283 20349
rect 2498 20340 2504 20352
rect 2556 20340 2562 20392
rect 2774 20380 2780 20392
rect 2735 20352 2780 20380
rect 2774 20340 2780 20352
rect 2832 20340 2838 20392
rect 26326 20380 26332 20392
rect 26287 20352 26332 20380
rect 26326 20340 26332 20352
rect 26384 20340 26390 20392
rect 26970 20340 26976 20392
rect 27028 20380 27034 20392
rect 27525 20383 27583 20389
rect 27525 20380 27537 20383
rect 27028 20352 27537 20380
rect 27028 20340 27034 20352
rect 27525 20349 27537 20352
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 30101 20383 30159 20389
rect 30101 20349 30113 20383
rect 30147 20380 30159 20383
rect 31496 20380 31524 20408
rect 30147 20352 31524 20380
rect 34885 20383 34943 20389
rect 30147 20349 30159 20352
rect 30101 20343 30159 20349
rect 34885 20349 34897 20383
rect 34931 20349 34943 20383
rect 35176 20380 35204 20411
rect 35802 20408 35808 20420
rect 35860 20408 35866 20460
rect 35989 20451 36047 20457
rect 35989 20417 36001 20451
rect 36035 20448 36047 20451
rect 36078 20448 36084 20460
rect 36035 20420 36084 20448
rect 36035 20417 36047 20420
rect 35989 20411 36047 20417
rect 36078 20408 36084 20420
rect 36136 20448 36142 20460
rect 36354 20448 36360 20460
rect 36136 20420 36360 20448
rect 36136 20408 36142 20420
rect 36354 20408 36360 20420
rect 36412 20408 36418 20460
rect 36449 20451 36507 20457
rect 36449 20417 36461 20451
rect 36495 20417 36507 20451
rect 36449 20411 36507 20417
rect 36262 20380 36268 20392
rect 35176 20352 36268 20380
rect 34885 20343 34943 20349
rect 34900 20312 34928 20343
rect 36262 20340 36268 20352
rect 36320 20380 36326 20392
rect 36464 20380 36492 20411
rect 37274 20408 37280 20460
rect 37332 20448 37338 20460
rect 38010 20457 38016 20460
rect 37737 20451 37795 20457
rect 37737 20448 37749 20451
rect 37332 20420 37749 20448
rect 37332 20408 37338 20420
rect 37737 20417 37749 20420
rect 37783 20417 37795 20451
rect 37737 20411 37795 20417
rect 38004 20411 38016 20457
rect 38068 20448 38074 20460
rect 40512 20457 40540 20488
rect 41598 20476 41604 20488
rect 41656 20476 41662 20528
rect 42536 20516 42564 20556
rect 42978 20544 42984 20556
rect 43036 20544 43042 20596
rect 42536 20488 43668 20516
rect 40497 20451 40555 20457
rect 38068 20420 38104 20448
rect 38010 20408 38016 20411
rect 38068 20408 38074 20420
rect 40497 20417 40509 20451
rect 40543 20417 40555 20451
rect 40497 20411 40555 20417
rect 40764 20451 40822 20457
rect 40764 20417 40776 20451
rect 40810 20448 40822 20451
rect 41322 20448 41328 20460
rect 40810 20420 41328 20448
rect 40810 20417 40822 20420
rect 40764 20411 40822 20417
rect 41322 20408 41328 20420
rect 41380 20408 41386 20460
rect 43257 20451 43315 20457
rect 43257 20417 43269 20451
rect 43303 20417 43315 20451
rect 43257 20411 43315 20417
rect 43349 20451 43407 20457
rect 43349 20417 43361 20451
rect 43395 20417 43407 20451
rect 43349 20411 43407 20417
rect 36320 20352 36492 20380
rect 36320 20340 36326 20352
rect 35897 20315 35955 20321
rect 35897 20312 35909 20315
rect 33244 20284 34376 20312
rect 34900 20284 35909 20312
rect 27522 20244 27528 20256
rect 27483 20216 27528 20244
rect 27522 20204 27528 20216
rect 27580 20204 27586 20256
rect 33042 20204 33048 20256
rect 33100 20244 33106 20256
rect 33244 20244 33272 20284
rect 33686 20244 33692 20256
rect 33100 20216 33272 20244
rect 33599 20216 33692 20244
rect 33100 20204 33106 20216
rect 33686 20204 33692 20216
rect 33744 20244 33750 20256
rect 34238 20244 34244 20256
rect 33744 20216 34244 20244
rect 33744 20204 33750 20216
rect 34238 20204 34244 20216
rect 34296 20204 34302 20256
rect 34348 20244 34376 20284
rect 35897 20281 35909 20284
rect 35943 20281 35955 20315
rect 40494 20312 40500 20324
rect 35897 20275 35955 20281
rect 38948 20284 40500 20312
rect 35986 20244 35992 20256
rect 34348 20216 35992 20244
rect 35986 20204 35992 20216
rect 36044 20204 36050 20256
rect 36538 20244 36544 20256
rect 36499 20216 36544 20244
rect 36538 20204 36544 20216
rect 36596 20204 36602 20256
rect 37734 20204 37740 20256
rect 37792 20244 37798 20256
rect 38102 20244 38108 20256
rect 37792 20216 38108 20244
rect 37792 20204 37798 20216
rect 38102 20204 38108 20216
rect 38160 20244 38166 20256
rect 38948 20244 38976 20284
rect 40494 20272 40500 20284
rect 40552 20272 40558 20324
rect 39114 20244 39120 20256
rect 38160 20216 38976 20244
rect 39075 20216 39120 20244
rect 38160 20204 38166 20216
rect 39114 20204 39120 20216
rect 39172 20204 39178 20256
rect 41874 20244 41880 20256
rect 41835 20216 41880 20244
rect 41874 20204 41880 20216
rect 41932 20204 41938 20256
rect 43272 20244 43300 20411
rect 43364 20324 43392 20411
rect 43438 20408 43444 20460
rect 43496 20448 43502 20460
rect 43640 20457 43668 20488
rect 43625 20451 43683 20457
rect 43496 20420 43541 20448
rect 43496 20408 43502 20420
rect 43625 20417 43637 20451
rect 43671 20417 43683 20451
rect 44082 20448 44088 20460
rect 44043 20420 44088 20448
rect 43625 20411 43683 20417
rect 44082 20408 44088 20420
rect 44140 20408 44146 20460
rect 44269 20451 44327 20457
rect 44269 20417 44281 20451
rect 44315 20448 44327 20451
rect 44634 20448 44640 20460
rect 44315 20420 44640 20448
rect 44315 20417 44327 20420
rect 44269 20411 44327 20417
rect 43346 20272 43352 20324
rect 43404 20272 43410 20324
rect 44284 20312 44312 20411
rect 44634 20408 44640 20420
rect 44692 20408 44698 20460
rect 47026 20448 47032 20460
rect 46987 20420 47032 20448
rect 47026 20408 47032 20420
rect 47084 20448 47090 20460
rect 47302 20448 47308 20460
rect 47084 20420 47308 20448
rect 47084 20408 47090 20420
rect 47302 20408 47308 20420
rect 47360 20408 47366 20460
rect 43456 20284 44312 20312
rect 43456 20244 43484 20284
rect 43272 20216 43484 20244
rect 43990 20204 43996 20256
rect 44048 20244 44054 20256
rect 44085 20247 44143 20253
rect 44085 20244 44097 20247
rect 44048 20216 44097 20244
rect 44048 20204 44054 20216
rect 44085 20213 44097 20216
rect 44131 20213 44143 20247
rect 44085 20207 44143 20213
rect 46658 20204 46664 20256
rect 46716 20244 46722 20256
rect 47121 20247 47179 20253
rect 47121 20244 47133 20247
rect 46716 20216 47133 20244
rect 46716 20204 46722 20216
rect 47121 20213 47133 20216
rect 47167 20213 47179 20247
rect 47946 20244 47952 20256
rect 47907 20216 47952 20244
rect 47121 20207 47179 20213
rect 47946 20204 47952 20216
rect 48004 20204 48010 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 2498 20040 2504 20052
rect 2459 20012 2504 20040
rect 2498 20000 2504 20012
rect 2556 20000 2562 20052
rect 32858 20040 32864 20052
rect 32819 20012 32864 20040
rect 32858 20000 32864 20012
rect 32916 20000 32922 20052
rect 33962 20000 33968 20052
rect 34020 20040 34026 20052
rect 34149 20043 34207 20049
rect 34149 20040 34161 20043
rect 34020 20012 34161 20040
rect 34020 20000 34026 20012
rect 34149 20009 34161 20012
rect 34195 20009 34207 20043
rect 34149 20003 34207 20009
rect 34333 20043 34391 20049
rect 34333 20009 34345 20043
rect 34379 20040 34391 20043
rect 34790 20040 34796 20052
rect 34379 20012 34796 20040
rect 34379 20009 34391 20012
rect 34333 20003 34391 20009
rect 34790 20000 34796 20012
rect 34848 20000 34854 20052
rect 34885 20043 34943 20049
rect 34885 20009 34897 20043
rect 34931 20040 34943 20043
rect 35802 20040 35808 20052
rect 34931 20012 35808 20040
rect 34931 20009 34943 20012
rect 34885 20003 34943 20009
rect 35802 20000 35808 20012
rect 35860 20000 35866 20052
rect 35894 20000 35900 20052
rect 35952 20040 35958 20052
rect 36170 20040 36176 20052
rect 35952 20012 36176 20040
rect 35952 20000 35958 20012
rect 36170 20000 36176 20012
rect 36228 20000 36234 20052
rect 37829 20043 37887 20049
rect 37829 20009 37841 20043
rect 37875 20040 37887 20043
rect 38010 20040 38016 20052
rect 37875 20012 38016 20040
rect 37875 20009 37887 20012
rect 37829 20003 37887 20009
rect 38010 20000 38016 20012
rect 38068 20000 38074 20052
rect 39022 20040 39028 20052
rect 38120 20012 38332 20040
rect 38983 20012 39028 20040
rect 34238 19932 34244 19984
rect 34296 19972 34302 19984
rect 34296 19944 36124 19972
rect 34296 19932 34302 19944
rect 33686 19904 33692 19916
rect 33152 19876 33692 19904
rect 2130 19796 2136 19848
rect 2188 19836 2194 19848
rect 2409 19839 2467 19845
rect 2409 19836 2421 19839
rect 2188 19808 2421 19836
rect 2188 19796 2194 19808
rect 2409 19805 2421 19808
rect 2455 19836 2467 19839
rect 3234 19836 3240 19848
rect 2455 19808 3240 19836
rect 2455 19805 2467 19808
rect 2409 19799 2467 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 33152 19845 33180 19876
rect 33686 19864 33692 19876
rect 33744 19864 33750 19916
rect 33137 19839 33195 19845
rect 33137 19805 33149 19839
rect 33183 19805 33195 19839
rect 33137 19799 33195 19805
rect 33229 19839 33287 19845
rect 33229 19805 33241 19839
rect 33275 19805 33287 19839
rect 33229 19799 33287 19805
rect 33244 19768 33272 19799
rect 33318 19796 33324 19848
rect 33376 19836 33382 19848
rect 33505 19839 33563 19845
rect 33376 19808 33421 19836
rect 33376 19796 33382 19808
rect 33505 19805 33517 19839
rect 33551 19836 33563 19839
rect 34606 19836 34612 19848
rect 33551 19808 34612 19836
rect 33551 19805 33563 19808
rect 33505 19799 33563 19805
rect 34606 19796 34612 19808
rect 34664 19796 34670 19848
rect 35069 19839 35127 19845
rect 35069 19836 35081 19839
rect 34900 19808 35081 19836
rect 33870 19768 33876 19780
rect 33244 19740 33876 19768
rect 33870 19728 33876 19740
rect 33928 19728 33934 19780
rect 33965 19771 34023 19777
rect 33965 19737 33977 19771
rect 34011 19768 34023 19771
rect 34330 19768 34336 19780
rect 34011 19740 34336 19768
rect 34011 19737 34023 19740
rect 33965 19731 34023 19737
rect 34330 19728 34336 19740
rect 34388 19768 34394 19780
rect 34698 19768 34704 19780
rect 34388 19740 34704 19768
rect 34388 19728 34394 19740
rect 34698 19728 34704 19740
rect 34756 19728 34762 19780
rect 34900 19768 34928 19808
rect 35069 19805 35081 19808
rect 35115 19805 35127 19839
rect 35069 19799 35127 19805
rect 35342 19796 35348 19848
rect 35400 19836 35406 19848
rect 35400 19808 35445 19836
rect 35400 19796 35406 19808
rect 35894 19796 35900 19848
rect 35952 19836 35958 19848
rect 35989 19839 36047 19845
rect 35989 19836 36001 19839
rect 35952 19808 36001 19836
rect 35952 19796 35958 19808
rect 35989 19805 36001 19808
rect 36035 19805 36047 19839
rect 36096 19836 36124 19944
rect 36262 19904 36268 19916
rect 36223 19876 36268 19904
rect 36262 19864 36268 19876
rect 36320 19864 36326 19916
rect 38120 19845 38148 20012
rect 38194 19932 38200 19984
rect 38252 19932 38258 19984
rect 38304 19972 38332 20012
rect 39022 20000 39028 20012
rect 39080 20000 39086 20052
rect 41322 20040 41328 20052
rect 41283 20012 41328 20040
rect 41322 20000 41328 20012
rect 41380 20000 41386 20052
rect 41966 20040 41972 20052
rect 41927 20012 41972 20040
rect 41966 20000 41972 20012
rect 42024 20000 42030 20052
rect 43257 20043 43315 20049
rect 43257 20009 43269 20043
rect 43303 20040 43315 20043
rect 43438 20040 43444 20052
rect 43303 20012 43444 20040
rect 43303 20009 43315 20012
rect 43257 20003 43315 20009
rect 43438 20000 43444 20012
rect 43496 20000 43502 20052
rect 38304 19944 38976 19972
rect 38212 19845 38240 19932
rect 38948 19904 38976 19944
rect 40126 19932 40132 19984
rect 40184 19972 40190 19984
rect 47946 19972 47952 19984
rect 40184 19944 43576 19972
rect 40184 19932 40190 19944
rect 39114 19904 39120 19916
rect 38948 19876 39120 19904
rect 36173 19839 36231 19845
rect 36173 19836 36185 19839
rect 36096 19808 36185 19836
rect 35989 19799 36047 19805
rect 36173 19805 36185 19808
rect 36219 19836 36231 19839
rect 36725 19839 36783 19845
rect 36725 19836 36737 19839
rect 36219 19808 36737 19836
rect 36219 19805 36231 19808
rect 36173 19799 36231 19805
rect 36725 19805 36737 19808
rect 36771 19805 36783 19839
rect 36725 19799 36783 19805
rect 38105 19839 38163 19845
rect 38105 19805 38117 19839
rect 38151 19805 38163 19839
rect 38105 19799 38163 19805
rect 38197 19839 38255 19845
rect 38197 19805 38209 19839
rect 38243 19805 38255 19839
rect 38197 19799 38255 19805
rect 38286 19796 38292 19848
rect 38344 19836 38350 19848
rect 38344 19808 38389 19836
rect 38344 19796 38350 19808
rect 38470 19796 38476 19848
rect 38528 19836 38534 19848
rect 38948 19845 38976 19876
rect 39114 19864 39120 19876
rect 39172 19904 39178 19916
rect 40405 19907 40463 19913
rect 40405 19904 40417 19907
rect 39172 19876 40417 19904
rect 39172 19864 39178 19876
rect 40405 19873 40417 19876
rect 40451 19873 40463 19907
rect 40405 19867 40463 19873
rect 40497 19907 40555 19913
rect 40497 19873 40509 19907
rect 40543 19904 40555 19907
rect 40543 19876 41920 19904
rect 40543 19873 40555 19876
rect 40497 19867 40555 19873
rect 41892 19848 41920 19876
rect 38933 19839 38991 19845
rect 38528 19808 38573 19836
rect 38528 19796 38534 19808
rect 38933 19805 38945 19839
rect 38979 19805 38991 19839
rect 38933 19799 38991 19805
rect 39482 19796 39488 19848
rect 39540 19836 39546 19848
rect 40126 19836 40132 19848
rect 39540 19808 40132 19836
rect 39540 19796 39546 19808
rect 40126 19796 40132 19808
rect 40184 19836 40190 19848
rect 40221 19839 40279 19845
rect 40221 19836 40233 19839
rect 40184 19808 40233 19836
rect 40184 19796 40190 19808
rect 40221 19805 40233 19808
rect 40267 19805 40279 19839
rect 41230 19836 41236 19848
rect 41191 19808 41236 19836
rect 40221 19799 40279 19805
rect 41230 19796 41236 19808
rect 41288 19796 41294 19848
rect 41322 19796 41328 19848
rect 41380 19836 41386 19848
rect 41874 19836 41880 19848
rect 41380 19808 41425 19836
rect 41835 19808 41880 19836
rect 41380 19796 41386 19808
rect 41874 19796 41880 19808
rect 41932 19796 41938 19848
rect 43162 19836 43168 19848
rect 43123 19808 43168 19836
rect 43162 19796 43168 19808
rect 43220 19796 43226 19848
rect 43346 19796 43352 19848
rect 43404 19836 43410 19848
rect 43548 19836 43576 19944
rect 46492 19944 47952 19972
rect 43809 19907 43867 19913
rect 43809 19873 43821 19907
rect 43855 19904 43867 19907
rect 44634 19904 44640 19916
rect 43855 19876 44640 19904
rect 43855 19873 43867 19876
rect 43809 19867 43867 19873
rect 44634 19864 44640 19876
rect 44692 19864 44698 19916
rect 46492 19913 46520 19944
rect 47946 19932 47952 19944
rect 48004 19932 48010 19984
rect 46477 19907 46535 19913
rect 46477 19873 46489 19907
rect 46523 19873 46535 19907
rect 46658 19904 46664 19916
rect 46619 19876 46664 19904
rect 46477 19867 46535 19873
rect 46658 19864 46664 19876
rect 46716 19864 46722 19916
rect 48222 19904 48228 19916
rect 48183 19876 48228 19904
rect 48222 19864 48228 19876
rect 48280 19864 48286 19916
rect 43993 19839 44051 19845
rect 43993 19836 44005 19839
rect 43404 19808 43497 19836
rect 43548 19808 44005 19836
rect 43404 19796 43410 19808
rect 43993 19805 44005 19808
rect 44039 19836 44051 19839
rect 44082 19836 44088 19848
rect 44039 19808 44088 19836
rect 44039 19805 44051 19808
rect 43993 19799 44051 19805
rect 44082 19796 44088 19808
rect 44140 19796 44146 19848
rect 34808 19740 34928 19768
rect 38580 19740 40264 19768
rect 34808 19712 34836 19740
rect 34175 19703 34233 19709
rect 34175 19669 34187 19703
rect 34221 19700 34233 19703
rect 34790 19700 34796 19712
rect 34221 19672 34796 19700
rect 34221 19669 34233 19672
rect 34175 19663 34233 19669
rect 34790 19660 34796 19672
rect 34848 19660 34854 19712
rect 34974 19660 34980 19712
rect 35032 19700 35038 19712
rect 35253 19703 35311 19709
rect 35253 19700 35265 19703
rect 35032 19672 35265 19700
rect 35032 19660 35038 19672
rect 35253 19669 35265 19672
rect 35299 19669 35311 19703
rect 35802 19700 35808 19712
rect 35763 19672 35808 19700
rect 35253 19663 35311 19669
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 36814 19700 36820 19712
rect 36775 19672 36820 19700
rect 36814 19660 36820 19672
rect 36872 19660 36878 19712
rect 38194 19660 38200 19712
rect 38252 19700 38258 19712
rect 38580 19700 38608 19740
rect 40034 19700 40040 19712
rect 38252 19672 38608 19700
rect 39995 19672 40040 19700
rect 38252 19660 38258 19672
rect 40034 19660 40040 19672
rect 40092 19660 40098 19712
rect 40236 19700 40264 19740
rect 40586 19728 40592 19780
rect 40644 19768 40650 19780
rect 40957 19771 41015 19777
rect 40957 19768 40969 19771
rect 40644 19740 40969 19768
rect 40644 19728 40650 19740
rect 40957 19737 40969 19740
rect 41003 19737 41015 19771
rect 43364 19768 43392 19796
rect 40957 19731 41015 19737
rect 41708 19740 43392 19768
rect 41708 19712 41736 19740
rect 41049 19703 41107 19709
rect 41049 19700 41061 19703
rect 40236 19672 41061 19700
rect 41049 19669 41061 19672
rect 41095 19700 41107 19703
rect 41690 19700 41696 19712
rect 41095 19672 41696 19700
rect 41095 19669 41107 19672
rect 41049 19663 41107 19669
rect 41690 19660 41696 19672
rect 41748 19660 41754 19712
rect 44177 19703 44235 19709
rect 44177 19669 44189 19703
rect 44223 19700 44235 19703
rect 44358 19700 44364 19712
rect 44223 19672 44364 19700
rect 44223 19669 44235 19672
rect 44177 19663 44235 19669
rect 44358 19660 44364 19672
rect 44416 19660 44422 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 33318 19456 33324 19508
rect 33376 19496 33382 19508
rect 34149 19499 34207 19505
rect 34149 19496 34161 19499
rect 33376 19468 34161 19496
rect 33376 19456 33382 19468
rect 34149 19465 34161 19468
rect 34195 19465 34207 19499
rect 35158 19496 35164 19508
rect 34149 19459 34207 19465
rect 34900 19468 35164 19496
rect 34900 19428 34928 19468
rect 35158 19456 35164 19468
rect 35216 19496 35222 19508
rect 35434 19496 35440 19508
rect 35216 19468 35440 19496
rect 35216 19456 35222 19468
rect 35434 19456 35440 19468
rect 35492 19496 35498 19508
rect 35492 19468 35940 19496
rect 35492 19456 35498 19468
rect 32876 19400 34928 19428
rect 32876 19369 32904 19400
rect 34974 19388 34980 19440
rect 35032 19428 35038 19440
rect 35710 19428 35716 19440
rect 35032 19400 35716 19428
rect 35032 19388 35038 19400
rect 32861 19363 32919 19369
rect 32861 19329 32873 19363
rect 32907 19329 32919 19363
rect 33042 19360 33048 19372
rect 33003 19332 33048 19360
rect 32861 19323 32919 19329
rect 33042 19320 33048 19332
rect 33100 19320 33106 19372
rect 35116 19369 35144 19400
rect 35710 19388 35716 19400
rect 35768 19388 35774 19440
rect 35912 19437 35940 19468
rect 36354 19456 36360 19508
rect 36412 19496 36418 19508
rect 37921 19499 37979 19505
rect 37921 19496 37933 19499
rect 36412 19468 37933 19496
rect 36412 19456 36418 19468
rect 37921 19465 37933 19468
rect 37967 19496 37979 19499
rect 38102 19496 38108 19508
rect 37967 19468 38108 19496
rect 37967 19465 37979 19468
rect 37921 19459 37979 19465
rect 38102 19456 38108 19468
rect 38160 19456 38166 19508
rect 38286 19456 38292 19508
rect 38344 19496 38350 19508
rect 38565 19499 38623 19505
rect 38565 19496 38577 19499
rect 38344 19468 38577 19496
rect 38344 19456 38350 19468
rect 38565 19465 38577 19468
rect 38611 19465 38623 19499
rect 38565 19459 38623 19465
rect 40129 19499 40187 19505
rect 40129 19465 40141 19499
rect 40175 19465 40187 19499
rect 41230 19496 41236 19508
rect 41191 19468 41236 19496
rect 40129 19459 40187 19465
rect 35897 19431 35955 19437
rect 35897 19397 35909 19431
rect 35943 19397 35955 19431
rect 35897 19391 35955 19397
rect 35986 19388 35992 19440
rect 36044 19428 36050 19440
rect 36081 19431 36139 19437
rect 36081 19428 36093 19431
rect 36044 19400 36093 19428
rect 36044 19388 36050 19400
rect 36081 19397 36093 19400
rect 36127 19397 36139 19431
rect 38746 19428 38752 19440
rect 36081 19391 36139 19397
rect 36372 19400 38752 19428
rect 33873 19363 33931 19369
rect 33152 19332 33824 19360
rect 32953 19295 33011 19301
rect 32953 19261 32965 19295
rect 32999 19292 33011 19295
rect 33152 19292 33180 19332
rect 33502 19292 33508 19304
rect 32999 19264 33180 19292
rect 33463 19264 33508 19292
rect 32999 19261 33011 19264
rect 32953 19255 33011 19261
rect 33502 19252 33508 19264
rect 33560 19252 33566 19304
rect 33796 19292 33824 19332
rect 33873 19329 33885 19363
rect 33919 19360 33931 19363
rect 35070 19363 35144 19369
rect 33919 19332 35020 19360
rect 33919 19329 33931 19332
rect 33873 19323 33931 19329
rect 33962 19292 33968 19304
rect 33796 19264 33968 19292
rect 33962 19252 33968 19264
rect 34020 19252 34026 19304
rect 34992 19224 35020 19332
rect 35070 19329 35082 19363
rect 35116 19332 35144 19363
rect 35345 19363 35403 19369
rect 35116 19329 35128 19332
rect 35070 19323 35128 19329
rect 35345 19329 35357 19363
rect 35391 19360 35403 19363
rect 35802 19360 35808 19372
rect 35391 19332 35808 19360
rect 35391 19329 35403 19332
rect 35345 19323 35403 19329
rect 35802 19320 35808 19332
rect 35860 19320 35866 19372
rect 35158 19292 35164 19304
rect 35119 19264 35164 19292
rect 35158 19252 35164 19264
rect 35216 19252 35222 19304
rect 35253 19295 35311 19301
rect 35253 19261 35265 19295
rect 35299 19292 35311 19295
rect 36004 19292 36032 19388
rect 35299 19264 36032 19292
rect 35299 19261 35311 19264
rect 35253 19255 35311 19261
rect 36265 19227 36323 19233
rect 36265 19224 36277 19227
rect 34992 19196 36277 19224
rect 36265 19193 36277 19196
rect 36311 19193 36323 19227
rect 36265 19187 36323 19193
rect 34885 19159 34943 19165
rect 34885 19125 34897 19159
rect 34931 19156 34943 19159
rect 36372 19156 36400 19400
rect 38746 19388 38752 19400
rect 38804 19428 38810 19440
rect 39942 19428 39948 19440
rect 38804 19400 39948 19428
rect 38804 19388 38810 19400
rect 39942 19388 39948 19400
rect 40000 19388 40006 19440
rect 40144 19428 40172 19459
rect 41230 19456 41236 19468
rect 41288 19456 41294 19508
rect 43162 19456 43168 19508
rect 43220 19496 43226 19508
rect 43717 19499 43775 19505
rect 43717 19496 43729 19499
rect 43220 19468 43729 19496
rect 43220 19456 43226 19468
rect 43717 19465 43729 19468
rect 43763 19465 43775 19499
rect 43717 19459 43775 19465
rect 43806 19456 43812 19508
rect 43864 19496 43870 19508
rect 44545 19499 44603 19505
rect 44545 19496 44557 19499
rect 43864 19468 44557 19496
rect 43864 19456 43870 19468
rect 44545 19465 44557 19468
rect 44591 19465 44603 19499
rect 44545 19459 44603 19465
rect 40144 19400 44680 19428
rect 38289 19363 38347 19369
rect 38289 19329 38301 19363
rect 38335 19360 38347 19363
rect 38930 19360 38936 19372
rect 38335 19332 38936 19360
rect 38335 19329 38347 19332
rect 38289 19323 38347 19329
rect 38930 19320 38936 19332
rect 38988 19320 38994 19372
rect 39025 19363 39083 19369
rect 39025 19329 39037 19363
rect 39071 19329 39083 19363
rect 39025 19323 39083 19329
rect 38381 19295 38439 19301
rect 38381 19261 38393 19295
rect 38427 19292 38439 19295
rect 38562 19292 38568 19304
rect 38427 19264 38568 19292
rect 38427 19261 38439 19264
rect 38381 19255 38439 19261
rect 38562 19252 38568 19264
rect 38620 19292 38626 19304
rect 39040 19292 39068 19323
rect 39114 19320 39120 19372
rect 39172 19360 39178 19372
rect 39393 19363 39451 19369
rect 39393 19360 39405 19363
rect 39172 19332 39405 19360
rect 39172 19320 39178 19332
rect 39393 19329 39405 19332
rect 39439 19329 39451 19363
rect 39393 19323 39451 19329
rect 39482 19320 39488 19372
rect 39540 19360 39546 19372
rect 39540 19332 39585 19360
rect 39540 19320 39546 19332
rect 40034 19320 40040 19372
rect 40092 19360 40098 19372
rect 40589 19363 40647 19369
rect 40589 19360 40601 19363
rect 40092 19332 40601 19360
rect 40092 19320 40098 19332
rect 40589 19329 40601 19332
rect 40635 19329 40647 19363
rect 40589 19323 40647 19329
rect 40678 19320 40684 19372
rect 40736 19360 40742 19372
rect 41141 19363 41199 19369
rect 41141 19360 41153 19363
rect 40736 19332 41153 19360
rect 40736 19320 40742 19332
rect 41141 19329 41153 19332
rect 41187 19329 41199 19363
rect 41141 19323 41199 19329
rect 41325 19363 41383 19369
rect 41325 19329 41337 19363
rect 41371 19360 41383 19363
rect 41874 19360 41880 19372
rect 41371 19332 41880 19360
rect 41371 19329 41383 19332
rect 41325 19323 41383 19329
rect 41874 19320 41880 19332
rect 41932 19320 41938 19372
rect 38620 19264 39068 19292
rect 38620 19252 38626 19264
rect 40218 19252 40224 19304
rect 40276 19292 40282 19304
rect 43272 19301 43300 19400
rect 43349 19363 43407 19369
rect 43349 19329 43361 19363
rect 43395 19360 43407 19363
rect 43806 19360 43812 19372
rect 43395 19332 43812 19360
rect 43395 19329 43407 19332
rect 43349 19323 43407 19329
rect 43806 19320 43812 19332
rect 43864 19320 43870 19372
rect 44358 19360 44364 19372
rect 44319 19332 44364 19360
rect 44358 19320 44364 19332
rect 44416 19320 44422 19372
rect 44652 19369 44680 19400
rect 44637 19363 44695 19369
rect 44637 19329 44649 19363
rect 44683 19329 44695 19363
rect 44637 19323 44695 19329
rect 47029 19363 47087 19369
rect 47029 19329 47041 19363
rect 47075 19360 47087 19363
rect 47210 19360 47216 19372
rect 47075 19332 47216 19360
rect 47075 19329 47087 19332
rect 47029 19323 47087 19329
rect 47210 19320 47216 19332
rect 47268 19360 47274 19372
rect 47670 19360 47676 19372
rect 47268 19332 47676 19360
rect 47268 19320 47274 19332
rect 47670 19320 47676 19332
rect 47728 19320 47734 19372
rect 40313 19295 40371 19301
rect 40313 19292 40325 19295
rect 40276 19264 40325 19292
rect 40276 19252 40282 19264
rect 40313 19261 40325 19264
rect 40359 19261 40371 19295
rect 40313 19255 40371 19261
rect 40405 19295 40463 19301
rect 40405 19261 40417 19295
rect 40451 19261 40463 19295
rect 40405 19255 40463 19261
rect 40497 19295 40555 19301
rect 40497 19261 40509 19295
rect 40543 19261 40555 19295
rect 40497 19255 40555 19261
rect 43257 19295 43315 19301
rect 43257 19261 43269 19295
rect 43303 19261 43315 19295
rect 43257 19255 43315 19261
rect 44177 19295 44235 19301
rect 44177 19261 44189 19295
rect 44223 19292 44235 19295
rect 44266 19292 44272 19304
rect 44223 19264 44272 19292
rect 44223 19261 44235 19264
rect 44177 19255 44235 19261
rect 38654 19184 38660 19236
rect 38712 19224 38718 19236
rect 40420 19224 40448 19255
rect 38712 19196 40448 19224
rect 38712 19184 38718 19196
rect 39666 19156 39672 19168
rect 34931 19128 36400 19156
rect 39627 19128 39672 19156
rect 34931 19125 34943 19128
rect 34885 19119 34943 19125
rect 39666 19116 39672 19128
rect 39724 19116 39730 19168
rect 39942 19116 39948 19168
rect 40000 19156 40006 19168
rect 40512 19156 40540 19255
rect 44266 19252 44272 19264
rect 44324 19252 44330 19304
rect 47118 19156 47124 19168
rect 40000 19128 40540 19156
rect 47079 19128 47124 19156
rect 40000 19116 40006 19128
rect 47118 19116 47124 19128
rect 47176 19116 47182 19168
rect 47946 19156 47952 19168
rect 47907 19128 47952 19156
rect 47946 19116 47952 19128
rect 48004 19116 48010 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 34241 18955 34299 18961
rect 34241 18921 34253 18955
rect 34287 18952 34299 18955
rect 34330 18952 34336 18964
rect 34287 18924 34336 18952
rect 34287 18921 34299 18924
rect 34241 18915 34299 18921
rect 34330 18912 34336 18924
rect 34388 18912 34394 18964
rect 35710 18952 35716 18964
rect 35671 18924 35716 18952
rect 35710 18912 35716 18924
rect 35768 18912 35774 18964
rect 38930 18952 38936 18964
rect 38891 18924 38936 18952
rect 38930 18912 38936 18924
rect 38988 18912 38994 18964
rect 43806 18952 43812 18964
rect 43767 18924 43812 18952
rect 43806 18912 43812 18924
rect 43864 18912 43870 18964
rect 39482 18884 39488 18896
rect 34164 18856 36216 18884
rect 2038 18708 2044 18760
rect 2096 18748 2102 18760
rect 34164 18757 34192 18856
rect 36188 18828 36216 18856
rect 37660 18856 39488 18884
rect 35529 18819 35587 18825
rect 35529 18785 35541 18819
rect 35575 18816 35587 18819
rect 35618 18816 35624 18828
rect 35575 18788 35624 18816
rect 35575 18785 35587 18788
rect 35529 18779 35587 18785
rect 35618 18776 35624 18788
rect 35676 18776 35682 18828
rect 36170 18776 36176 18828
rect 36228 18816 36234 18828
rect 37660 18825 37688 18856
rect 39482 18844 39488 18856
rect 39540 18844 39546 18896
rect 40586 18884 40592 18896
rect 40547 18856 40592 18884
rect 40586 18844 40592 18856
rect 40644 18844 40650 18896
rect 47946 18884 47952 18896
rect 46492 18856 47952 18884
rect 37645 18819 37703 18825
rect 37645 18816 37657 18819
rect 36228 18788 37657 18816
rect 36228 18776 36234 18788
rect 37645 18785 37657 18788
rect 37691 18785 37703 18819
rect 39022 18816 39028 18828
rect 37645 18779 37703 18785
rect 37752 18788 39028 18816
rect 2317 18751 2375 18757
rect 2317 18748 2329 18751
rect 2096 18720 2329 18748
rect 2096 18708 2102 18720
rect 2317 18717 2329 18720
rect 2363 18717 2375 18751
rect 2317 18711 2375 18717
rect 34149 18751 34207 18757
rect 34149 18717 34161 18751
rect 34195 18717 34207 18751
rect 34149 18711 34207 18717
rect 34238 18708 34244 18760
rect 34296 18748 34302 18760
rect 34333 18751 34391 18757
rect 34333 18748 34345 18751
rect 34296 18720 34345 18748
rect 34296 18708 34302 18720
rect 34333 18717 34345 18720
rect 34379 18717 34391 18751
rect 34333 18711 34391 18717
rect 35437 18751 35495 18757
rect 35437 18717 35449 18751
rect 35483 18748 35495 18751
rect 36538 18748 36544 18760
rect 35483 18720 36544 18748
rect 35483 18717 35495 18720
rect 35437 18711 35495 18717
rect 36538 18708 36544 18720
rect 36596 18708 36602 18760
rect 37752 18757 37780 18788
rect 39022 18776 39028 18788
rect 39080 18776 39086 18828
rect 39666 18776 39672 18828
rect 39724 18816 39730 18828
rect 40129 18819 40187 18825
rect 40129 18816 40141 18819
rect 39724 18788 40141 18816
rect 39724 18776 39730 18788
rect 40129 18785 40141 18788
rect 40175 18785 40187 18819
rect 44358 18816 44364 18828
rect 40129 18779 40187 18785
rect 43824 18788 44364 18816
rect 37737 18751 37795 18757
rect 37737 18717 37749 18751
rect 37783 18717 37795 18751
rect 37737 18711 37795 18717
rect 38565 18751 38623 18757
rect 38565 18717 38577 18751
rect 38611 18748 38623 18751
rect 38654 18748 38660 18760
rect 38611 18720 38660 18748
rect 38611 18717 38623 18720
rect 38565 18711 38623 18717
rect 38105 18615 38163 18621
rect 38105 18581 38117 18615
rect 38151 18612 38163 18615
rect 38580 18612 38608 18711
rect 38654 18708 38660 18720
rect 38712 18708 38718 18760
rect 38746 18708 38752 18760
rect 38804 18748 38810 18760
rect 40218 18748 40224 18760
rect 38804 18720 38849 18748
rect 40179 18720 40224 18748
rect 38804 18708 38810 18720
rect 40218 18708 40224 18720
rect 40276 18708 40282 18760
rect 43824 18757 43852 18788
rect 44358 18776 44364 18788
rect 44416 18776 44422 18828
rect 46492 18825 46520 18856
rect 47946 18844 47952 18856
rect 48004 18844 48010 18896
rect 46477 18819 46535 18825
rect 46477 18785 46489 18819
rect 46523 18785 46535 18819
rect 46477 18779 46535 18785
rect 46661 18819 46719 18825
rect 46661 18785 46673 18819
rect 46707 18816 46719 18819
rect 47118 18816 47124 18828
rect 46707 18788 47124 18816
rect 46707 18785 46719 18788
rect 46661 18779 46719 18785
rect 47118 18776 47124 18788
rect 47176 18776 47182 18828
rect 48222 18816 48228 18828
rect 48183 18788 48228 18816
rect 48222 18776 48228 18788
rect 48280 18776 48286 18828
rect 43809 18751 43867 18757
rect 43809 18717 43821 18751
rect 43855 18717 43867 18751
rect 43990 18748 43996 18760
rect 43951 18720 43996 18748
rect 43809 18711 43867 18717
rect 43990 18708 43996 18720
rect 44048 18708 44054 18760
rect 38151 18584 38608 18612
rect 38151 18581 38163 18584
rect 38105 18575 38163 18581
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 35434 18408 35440 18420
rect 35395 18380 35440 18408
rect 35434 18368 35440 18380
rect 35492 18368 35498 18420
rect 38562 18408 38568 18420
rect 38523 18380 38568 18408
rect 38562 18368 38568 18380
rect 38620 18368 38626 18420
rect 38654 18368 38660 18420
rect 38712 18368 38718 18420
rect 40218 18368 40224 18420
rect 40276 18408 40282 18420
rect 40405 18411 40463 18417
rect 40405 18408 40417 18411
rect 40276 18380 40417 18408
rect 40276 18368 40282 18380
rect 40405 18377 40417 18380
rect 40451 18377 40463 18411
rect 40405 18371 40463 18377
rect 38672 18340 38700 18368
rect 38488 18312 38700 18340
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 35069 18275 35127 18281
rect 35069 18241 35081 18275
rect 35115 18272 35127 18275
rect 36814 18272 36820 18284
rect 35115 18244 36820 18272
rect 35115 18241 35127 18244
rect 35069 18235 35127 18241
rect 36814 18232 36820 18244
rect 36872 18232 36878 18284
rect 38488 18281 38516 18312
rect 38473 18275 38531 18281
rect 38473 18241 38485 18275
rect 38519 18241 38531 18275
rect 38473 18235 38531 18241
rect 38657 18275 38715 18281
rect 38657 18241 38669 18275
rect 38703 18272 38715 18275
rect 38746 18272 38752 18284
rect 38703 18244 38752 18272
rect 38703 18241 38715 18244
rect 38657 18235 38715 18241
rect 38746 18232 38752 18244
rect 38804 18232 38810 18284
rect 40037 18275 40095 18281
rect 40037 18241 40049 18275
rect 40083 18272 40095 18275
rect 41966 18272 41972 18284
rect 40083 18244 41972 18272
rect 40083 18241 40095 18244
rect 40037 18235 40095 18241
rect 41966 18232 41972 18244
rect 42024 18232 42030 18284
rect 47486 18232 47492 18284
rect 47544 18272 47550 18284
rect 47765 18275 47823 18281
rect 47765 18272 47777 18275
rect 47544 18244 47777 18272
rect 47544 18232 47550 18244
rect 47765 18241 47777 18244
rect 47811 18241 47823 18275
rect 47765 18235 47823 18241
rect 2222 18204 2228 18216
rect 2183 18176 2228 18204
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 2774 18204 2780 18216
rect 2735 18176 2780 18204
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 35161 18207 35219 18213
rect 35161 18173 35173 18207
rect 35207 18204 35219 18207
rect 35618 18204 35624 18216
rect 35207 18176 35624 18204
rect 35207 18173 35219 18176
rect 35161 18167 35219 18173
rect 35618 18164 35624 18176
rect 35676 18164 35682 18216
rect 40126 18204 40132 18216
rect 40087 18176 40132 18204
rect 40126 18164 40132 18176
rect 40184 18164 40190 18216
rect 47854 18068 47860 18080
rect 47815 18040 47860 18068
rect 47854 18028 47860 18040
rect 47912 18028 47918 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 2685 17867 2743 17873
rect 2685 17864 2697 17867
rect 2280 17836 2697 17864
rect 2280 17824 2286 17836
rect 2685 17833 2697 17836
rect 2731 17833 2743 17867
rect 2685 17827 2743 17833
rect 46661 17731 46719 17737
rect 46661 17697 46673 17731
rect 46707 17728 46719 17731
rect 47854 17728 47860 17740
rect 46707 17700 47860 17728
rect 46707 17697 46719 17700
rect 46661 17691 46719 17697
rect 47854 17688 47860 17700
rect 47912 17688 47918 17740
rect 48222 17728 48228 17740
rect 48183 17700 48228 17728
rect 48222 17688 48228 17700
rect 48280 17688 48286 17740
rect 2498 17620 2504 17672
rect 2556 17660 2562 17672
rect 2593 17663 2651 17669
rect 2593 17660 2605 17663
rect 2556 17632 2605 17660
rect 2556 17620 2562 17632
rect 2593 17629 2605 17632
rect 2639 17660 2651 17663
rect 4614 17660 4620 17672
rect 2639 17632 4620 17660
rect 2639 17629 2651 17632
rect 2593 17623 2651 17629
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 46474 17660 46480 17672
rect 46435 17632 46480 17660
rect 46474 17620 46480 17632
rect 46532 17620 46538 17672
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 2225 17255 2283 17261
rect 2225 17221 2237 17255
rect 2271 17252 2283 17255
rect 2866 17252 2872 17264
rect 2271 17224 2872 17252
rect 2271 17221 2283 17224
rect 2225 17215 2283 17221
rect 2866 17212 2872 17224
rect 2924 17212 2930 17264
rect 46474 17144 46480 17196
rect 46532 17184 46538 17196
rect 47949 17187 48007 17193
rect 47949 17184 47961 17187
rect 46532 17156 47961 17184
rect 46532 17144 46538 17156
rect 47949 17153 47961 17156
rect 47995 17153 48007 17187
rect 47949 17147 48007 17153
rect 2038 17116 2044 17128
rect 1999 17088 2044 17116
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 46474 16940 46480 16992
rect 46532 16980 46538 16992
rect 47213 16983 47271 16989
rect 47213 16980 47225 16983
rect 46532 16952 47225 16980
rect 46532 16940 46538 16952
rect 47213 16949 47225 16952
rect 47259 16949 47271 16983
rect 47213 16943 47271 16949
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 2317 16779 2375 16785
rect 2317 16776 2329 16779
rect 2096 16748 2329 16776
rect 2096 16736 2102 16748
rect 2317 16745 2329 16748
rect 2363 16745 2375 16779
rect 2317 16739 2375 16745
rect 2590 16600 2596 16652
rect 2648 16640 2654 16652
rect 3786 16640 3792 16652
rect 2648 16612 3792 16640
rect 2648 16600 2654 16612
rect 2792 16581 2820 16612
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 46474 16640 46480 16652
rect 46435 16612 46480 16640
rect 46474 16600 46480 16612
rect 46532 16600 46538 16652
rect 48222 16640 48228 16652
rect 48183 16612 48228 16640
rect 48222 16600 48228 16612
rect 48280 16600 48286 16652
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16574 2835 16575
rect 2823 16546 2857 16574
rect 2823 16541 2835 16546
rect 2777 16535 2835 16541
rect 2866 16504 2872 16516
rect 2827 16476 2872 16504
rect 2866 16464 2872 16476
rect 2924 16464 2930 16516
rect 46661 16507 46719 16513
rect 46661 16473 46673 16507
rect 46707 16504 46719 16507
rect 47854 16504 47860 16516
rect 46707 16476 47860 16504
rect 46707 16473 46719 16476
rect 46661 16467 46719 16473
rect 47854 16464 47860 16476
rect 47912 16464 47918 16516
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 47854 16232 47860 16244
rect 47815 16204 47860 16232
rect 47854 16192 47860 16204
rect 47912 16192 47918 16244
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1946 15484 1952 15496
rect 1907 15456 1952 15484
rect 1946 15444 1952 15456
rect 2004 15444 2010 15496
rect 2130 15444 2136 15496
rect 2188 15484 2194 15496
rect 2409 15487 2467 15493
rect 2409 15484 2421 15487
rect 2188 15456 2421 15484
rect 2188 15444 2194 15456
rect 2409 15453 2421 15456
rect 2455 15484 2467 15487
rect 2590 15484 2596 15496
rect 2455 15456 2596 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 47670 15484 47676 15496
rect 47631 15456 47676 15484
rect 47670 15444 47676 15456
rect 47728 15444 47734 15496
rect 2222 15308 2228 15360
rect 2280 15348 2286 15360
rect 2501 15351 2559 15357
rect 2501 15348 2513 15351
rect 2280 15320 2513 15348
rect 2280 15308 2286 15320
rect 2501 15317 2513 15320
rect 2547 15317 2559 15351
rect 2501 15311 2559 15317
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 2222 15076 2228 15088
rect 2183 15048 2228 15076
rect 2222 15036 2228 15048
rect 2280 15036 2286 15088
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 2004 14980 2053 15008
rect 2004 14968 2010 14980
rect 2041 14977 2053 14980
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 47486 14968 47492 15020
rect 47544 15008 47550 15020
rect 47765 15011 47823 15017
rect 47765 15008 47777 15011
rect 47544 14980 47777 15008
rect 47544 14968 47550 14980
rect 47765 14977 47777 14980
rect 47811 14977 47823 15011
rect 47765 14971 47823 14977
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 46658 14764 46664 14816
rect 46716 14804 46722 14816
rect 47857 14807 47915 14813
rect 47857 14804 47869 14807
rect 46716 14776 47869 14804
rect 46716 14764 46722 14776
rect 47857 14773 47869 14776
rect 47903 14773 47915 14807
rect 47857 14767 47915 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 47670 14532 47676 14544
rect 46492 14504 47676 14532
rect 2774 14464 2780 14476
rect 2735 14436 2780 14464
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 46492 14473 46520 14504
rect 47670 14492 47676 14504
rect 47728 14492 47734 14544
rect 46477 14467 46535 14473
rect 46477 14433 46489 14467
rect 46523 14433 46535 14467
rect 46658 14464 46664 14476
rect 46619 14436 46664 14464
rect 46477 14427 46535 14433
rect 46658 14424 46664 14436
rect 46716 14424 46722 14476
rect 48222 14464 48228 14476
rect 48183 14436 48228 14464
rect 48222 14424 48228 14436
rect 48280 14424 48286 14476
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 1762 14328 1768 14340
rect 1723 14300 1768 14328
rect 1762 14288 1768 14300
rect 1820 14288 1826 14340
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1762 14016 1768 14068
rect 1820 14056 1826 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 1820 14028 2881 14056
rect 1820 14016 1826 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 2317 13923 2375 13929
rect 2317 13920 2329 13923
rect 1636 13892 2329 13920
rect 1636 13880 1642 13892
rect 2317 13889 2329 13892
rect 2363 13889 2375 13923
rect 2317 13883 2375 13889
rect 2682 13880 2688 13932
rect 2740 13920 2746 13932
rect 2777 13923 2835 13929
rect 2777 13920 2789 13923
rect 2740 13892 2789 13920
rect 2740 13880 2746 13892
rect 2777 13889 2789 13892
rect 2823 13920 2835 13923
rect 3050 13920 3056 13932
rect 2823 13892 3056 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 47029 13923 47087 13929
rect 47029 13889 47041 13923
rect 47075 13920 47087 13923
rect 47486 13920 47492 13932
rect 47075 13892 47492 13920
rect 47075 13889 47087 13892
rect 47029 13883 47087 13889
rect 47486 13880 47492 13892
rect 47544 13880 47550 13932
rect 47118 13716 47124 13728
rect 47079 13688 47124 13716
rect 47118 13676 47124 13688
rect 47176 13676 47182 13728
rect 47946 13716 47952 13728
rect 47907 13688 47952 13716
rect 47946 13676 47952 13688
rect 48004 13676 48010 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 47946 13444 47952 13456
rect 46492 13416 47952 13444
rect 46492 13385 46520 13416
rect 47946 13404 47952 13416
rect 48004 13404 48010 13456
rect 46477 13379 46535 13385
rect 46477 13345 46489 13379
rect 46523 13345 46535 13379
rect 46477 13339 46535 13345
rect 46661 13379 46719 13385
rect 46661 13345 46673 13379
rect 46707 13376 46719 13379
rect 47118 13376 47124 13388
rect 46707 13348 47124 13376
rect 46707 13345 46719 13348
rect 46661 13339 46719 13345
rect 47118 13336 47124 13348
rect 47176 13336 47182 13388
rect 48222 13376 48228 13388
rect 48183 13348 48228 13376
rect 48222 13336 48228 13348
rect 48280 13336 48286 13388
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 46934 12792 46940 12844
rect 46992 12832 46998 12844
rect 47029 12835 47087 12841
rect 47029 12832 47041 12835
rect 46992 12804 47041 12832
rect 46992 12792 46998 12804
rect 47029 12801 47041 12804
rect 47075 12801 47087 12835
rect 47029 12795 47087 12801
rect 47118 12628 47124 12640
rect 47079 12600 47124 12628
rect 47118 12588 47124 12600
rect 47176 12588 47182 12640
rect 47946 12628 47952 12640
rect 47907 12600 47952 12628
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 47946 12356 47952 12368
rect 46492 12328 47952 12356
rect 46492 12297 46520 12328
rect 47946 12316 47952 12328
rect 48004 12316 48010 12368
rect 46477 12291 46535 12297
rect 46477 12257 46489 12291
rect 46523 12257 46535 12291
rect 46477 12251 46535 12257
rect 46661 12291 46719 12297
rect 46661 12257 46673 12291
rect 46707 12288 46719 12291
rect 47118 12288 47124 12300
rect 46707 12260 47124 12288
rect 46707 12257 46719 12260
rect 46661 12251 46719 12257
rect 47118 12248 47124 12260
rect 47176 12248 47182 12300
rect 48222 12288 48228 12300
rect 48183 12260 48228 12288
rect 48222 12248 48228 12260
rect 48280 12248 48286 12300
rect 2314 12220 2320 12232
rect 2275 12192 2320 12220
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 2314 11812 2320 11824
rect 2056 11784 2320 11812
rect 2056 11753 2084 11784
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11713 2099 11747
rect 47026 11744 47032 11756
rect 46987 11716 47032 11744
rect 2041 11707 2099 11713
rect 47026 11704 47032 11716
rect 47084 11704 47090 11756
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11676 2283 11679
rect 2314 11676 2320 11688
rect 2271 11648 2320 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 2832 11648 2877 11676
rect 2832 11636 2838 11648
rect 46658 11500 46664 11552
rect 46716 11540 46722 11552
rect 47121 11543 47179 11549
rect 47121 11540 47133 11543
rect 46716 11512 47133 11540
rect 46716 11500 46722 11512
rect 47121 11509 47133 11512
rect 47167 11509 47179 11543
rect 47946 11540 47952 11552
rect 47907 11512 47952 11540
rect 47121 11503 47179 11509
rect 47946 11500 47952 11512
rect 48004 11500 48010 11552
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 47946 11268 47952 11280
rect 46492 11240 47952 11268
rect 46492 11209 46520 11240
rect 47946 11228 47952 11240
rect 48004 11228 48010 11280
rect 46477 11203 46535 11209
rect 46477 11169 46489 11203
rect 46523 11169 46535 11203
rect 46658 11200 46664 11212
rect 46619 11172 46664 11200
rect 46477 11163 46535 11169
rect 46658 11160 46664 11172
rect 46716 11160 46722 11212
rect 46842 11160 46848 11212
rect 46900 11200 46906 11212
rect 46937 11203 46995 11209
rect 46937 11200 46949 11203
rect 46900 11172 46949 11200
rect 46900 11160 46906 11172
rect 46937 11169 46949 11172
rect 46983 11169 46995 11203
rect 46937 11163 46995 11169
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2958 11132 2964 11144
rect 2271 11104 2964 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 2188 10016 2329 10044
rect 2188 10004 2194 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3142 10044 3148 10056
rect 2823 10016 3148 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3142 10004 3148 10016
rect 3200 10044 3206 10056
rect 41414 10044 41420 10056
rect 3200 10016 41420 10044
rect 3200 10004 3206 10016
rect 41414 10004 41420 10016
rect 41472 10004 41478 10056
rect 2866 9908 2872 9920
rect 2827 9880 2872 9908
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 2317 9639 2375 9645
rect 2317 9605 2329 9639
rect 2363 9636 2375 9639
rect 2866 9636 2872 9648
rect 2363 9608 2872 9636
rect 2363 9605 2375 9608
rect 2317 9599 2375 9605
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 41414 9596 41420 9648
rect 41472 9636 41478 9648
rect 45186 9636 45192 9648
rect 41472 9608 45192 9636
rect 41472 9596 41478 9608
rect 45186 9596 45192 9608
rect 45244 9636 45250 9648
rect 47762 9636 47768 9648
rect 45244 9608 47768 9636
rect 45244 9596 45250 9608
rect 47762 9596 47768 9608
rect 47820 9596 47826 9648
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 2130 8956 2136 8968
rect 2091 8928 2136 8956
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2498 8916 2504 8968
rect 2556 8956 2562 8968
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 2556 8928 2605 8956
rect 2556 8916 2562 8928
rect 2593 8925 2605 8928
rect 2639 8956 2651 8959
rect 4614 8956 4620 8968
rect 2639 8928 4620 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2372 8792 2697 8820
rect 2372 8780 2378 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2685 8783 2743 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 2314 8548 2320 8560
rect 2275 8520 2320 8548
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 41233 8483 41291 8489
rect 41233 8449 41245 8483
rect 41279 8480 41291 8483
rect 44358 8480 44364 8492
rect 41279 8452 44364 8480
rect 41279 8449 41291 8452
rect 41233 8443 41291 8449
rect 44358 8440 44364 8452
rect 44416 8440 44422 8492
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 41414 8412 41420 8424
rect 2832 8384 2877 8412
rect 41375 8384 41420 8412
rect 2832 8372 2838 8384
rect 41414 8372 41420 8384
rect 41472 8372 41478 8424
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 4065 8007 4123 8013
rect 4065 8004 4077 8007
rect 2746 7976 4077 8004
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2746 7936 2774 7976
rect 4065 7973 4077 7976
rect 4111 7973 4123 8007
rect 4065 7967 4123 7973
rect 2958 7936 2964 7948
rect 1811 7908 2774 7936
rect 2919 7908 2964 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 47486 7936 47492 7948
rect 47447 7908 47492 7936
rect 47486 7896 47492 7908
rect 47544 7896 47550 7948
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 5810 7868 5816 7880
rect 4019 7840 5816 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 3988 7800 4016 7831
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 46014 7828 46020 7880
rect 46072 7868 46078 7880
rect 47765 7871 47823 7877
rect 47765 7868 47777 7871
rect 46072 7840 47777 7868
rect 46072 7828 46078 7840
rect 47765 7837 47777 7840
rect 47811 7837 47823 7871
rect 47765 7831 47823 7837
rect 2464 7772 4016 7800
rect 2464 7760 2470 7772
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 2225 7463 2283 7469
rect 2225 7429 2237 7463
rect 2271 7460 2283 7463
rect 4062 7460 4068 7472
rect 2271 7432 4068 7460
rect 2271 7429 2283 7432
rect 2225 7423 2283 7429
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4614 7392 4620 7404
rect 4571 7364 4620 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4614 7352 4620 7364
rect 4672 7392 4678 7404
rect 24578 7392 24584 7404
rect 4672 7364 24584 7392
rect 4672 7352 4678 7364
rect 24578 7352 24584 7364
rect 24636 7352 24642 7404
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 2056 7256 2084 7287
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 5074 7324 5080 7336
rect 2832 7296 2877 7324
rect 5035 7296 5080 7324
rect 2832 7284 2838 7296
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 2958 7256 2964 7268
rect 2056 7228 2964 7256
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 5074 7188 5080 7200
rect 1728 7160 5080 7188
rect 1728 7148 1734 7160
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 47946 7188 47952 7200
rect 47907 7160 47952 7188
rect 47946 7148 47952 7160
rect 48004 7148 48010 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 2317 6987 2375 6993
rect 2317 6984 2329 6987
rect 1636 6956 2329 6984
rect 1636 6944 1642 6956
rect 2317 6953 2329 6956
rect 2363 6953 2375 6987
rect 2317 6947 2375 6953
rect 47946 6916 47952 6928
rect 46860 6888 47952 6916
rect 2958 6848 2964 6860
rect 2919 6820 2964 6848
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 46477 6851 46535 6857
rect 46477 6817 46489 6851
rect 46523 6848 46535 6851
rect 46860 6848 46888 6888
rect 47946 6876 47952 6888
rect 48004 6876 48010 6928
rect 48222 6848 48228 6860
rect 46523 6820 46888 6848
rect 48183 6820 48228 6848
rect 46523 6817 46535 6820
rect 46477 6811 46535 6817
rect 48222 6808 48228 6820
rect 48280 6808 48286 6860
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3970 6780 3976 6792
rect 3108 6752 3976 6780
rect 3108 6740 3114 6752
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 46661 6715 46719 6721
rect 46661 6681 46673 6715
rect 46707 6712 46719 6715
rect 47854 6712 47860 6724
rect 46707 6684 47860 6712
rect 46707 6681 46719 6684
rect 46661 6675 46719 6681
rect 47854 6672 47860 6684
rect 47912 6672 47918 6724
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 47854 6440 47860 6452
rect 47815 6412 47860 6440
rect 47854 6400 47860 6412
rect 47912 6400 47918 6452
rect 47578 6372 47584 6384
rect 46400 6344 47584 6372
rect 46400 6313 46428 6344
rect 47578 6332 47584 6344
rect 47636 6332 47642 6384
rect 46385 6307 46443 6313
rect 46385 6273 46397 6307
rect 46431 6273 46443 6307
rect 46385 6267 46443 6273
rect 47029 6307 47087 6313
rect 47029 6273 47041 6307
rect 47075 6304 47087 6307
rect 47210 6304 47216 6316
rect 47075 6276 47216 6304
rect 47075 6273 47087 6276
rect 47029 6267 47087 6273
rect 47210 6264 47216 6276
rect 47268 6264 47274 6316
rect 47394 6264 47400 6316
rect 47452 6304 47458 6316
rect 47765 6307 47823 6313
rect 47765 6304 47777 6307
rect 47452 6276 47777 6304
rect 47452 6264 47458 6276
rect 47765 6273 47777 6276
rect 47811 6304 47823 6307
rect 48038 6304 48044 6316
rect 47811 6276 48044 6304
rect 47811 6273 47823 6276
rect 47765 6267 47823 6273
rect 48038 6264 48044 6276
rect 48096 6264 48102 6316
rect 2130 6236 2136 6248
rect 2091 6208 2136 6236
rect 2130 6196 2136 6208
rect 2188 6196 2194 6248
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 2866 6236 2872 6248
rect 2363 6208 2872 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3016 6208 3061 6236
rect 3016 6196 3022 6208
rect 4617 6103 4675 6109
rect 4617 6069 4629 6103
rect 4663 6100 4675 6103
rect 4982 6100 4988 6112
rect 4663 6072 4988 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 46474 6100 46480 6112
rect 46435 6072 46480 6100
rect 46474 6060 46480 6072
rect 46532 6060 46538 6112
rect 46658 6060 46664 6112
rect 46716 6100 46722 6112
rect 47121 6103 47179 6109
rect 47121 6100 47133 6103
rect 46716 6072 47133 6100
rect 46716 6060 46722 6072
rect 47121 6069 47133 6072
rect 47167 6069 47179 6103
rect 47121 6063 47179 6069
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 2188 5868 2329 5896
rect 2188 5856 2194 5868
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 2866 5896 2872 5908
rect 2827 5868 2872 5896
rect 2317 5859 2375 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 4028 5800 12434 5828
rect 4028 5788 4034 5800
rect 3988 5760 4016 5788
rect 2792 5732 4016 5760
rect 2792 5701 2820 5732
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 5445 5763 5503 5769
rect 5445 5760 5457 5763
rect 4764 5732 5457 5760
rect 4764 5720 4770 5732
rect 5445 5729 5457 5732
rect 5491 5729 5503 5763
rect 12406 5760 12434 5800
rect 17402 5760 17408 5772
rect 12406 5732 17408 5760
rect 5445 5723 5503 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 46658 5760 46664 5772
rect 46619 5732 46664 5760
rect 46658 5720 46664 5732
rect 46716 5720 46722 5772
rect 48222 5760 48228 5772
rect 48183 5732 48228 5760
rect 48222 5720 48228 5732
rect 48280 5720 48286 5772
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3844 5664 3985 5692
rect 3844 5652 3850 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 4798 5692 4804 5704
rect 4759 5664 4804 5692
rect 3973 5655 4031 5661
rect 3988 5624 4016 5655
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 46014 5692 46020 5704
rect 45975 5664 46020 5692
rect 46014 5652 46020 5664
rect 46072 5652 46078 5704
rect 46477 5695 46535 5701
rect 46477 5661 46489 5695
rect 46523 5661 46535 5695
rect 46477 5655 46535 5661
rect 10410 5624 10416 5636
rect 3988 5596 10416 5624
rect 10410 5584 10416 5596
rect 10468 5584 10474 5636
rect 46492 5624 46520 5655
rect 47946 5624 47952 5636
rect 46492 5596 47952 5624
rect 47946 5584 47952 5596
rect 48004 5584 48010 5636
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 4798 5352 4804 5364
rect 2148 5324 4804 5352
rect 2148 5225 2176 5324
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 2317 5287 2375 5293
rect 2317 5253 2329 5287
rect 2363 5284 2375 5287
rect 4062 5284 4068 5296
rect 2363 5256 4068 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 46014 5284 46020 5296
rect 45388 5256 46020 5284
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5718 5216 5724 5228
rect 5215 5188 5724 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 4448 5148 4476 5179
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 45388 5225 45416 5256
rect 46014 5244 46020 5256
rect 46072 5244 46078 5296
rect 45373 5219 45431 5225
rect 5868 5188 5913 5216
rect 5868 5176 5874 5188
rect 45373 5185 45385 5219
rect 45419 5185 45431 5219
rect 47946 5216 47952 5228
rect 47907 5188 47952 5216
rect 45373 5179 45431 5185
rect 47946 5176 47952 5188
rect 48004 5176 48010 5228
rect 5074 5148 5080 5160
rect 2832 5120 2877 5148
rect 4448 5120 5080 5148
rect 2832 5108 2838 5120
rect 5074 5108 5080 5120
rect 5132 5148 5138 5160
rect 8294 5148 8300 5160
rect 5132 5120 8300 5148
rect 5132 5108 5138 5120
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 44542 5108 44548 5160
rect 44600 5148 44606 5160
rect 45557 5151 45615 5157
rect 45557 5148 45569 5151
rect 44600 5120 45569 5148
rect 44600 5108 44606 5120
rect 45557 5117 45569 5120
rect 45603 5117 45615 5151
rect 45557 5111 45615 5117
rect 47213 5151 47271 5157
rect 47213 5117 47225 5151
rect 47259 5148 47271 5151
rect 48958 5148 48964 5160
rect 47259 5120 48964 5148
rect 47259 5117 47271 5120
rect 47213 5111 47271 5117
rect 48958 5108 48964 5120
rect 49016 5108 49022 5160
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 4798 5012 4804 5024
rect 4571 4984 4804 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 4948 4984 5273 5012
rect 4948 4972 4954 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 5261 4975 5319 4981
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5905 5015 5963 5021
rect 5905 5012 5917 5015
rect 5684 4984 5917 5012
rect 5684 4972 5690 4984
rect 5905 4981 5917 4984
rect 5951 4981 5963 5015
rect 5905 4975 5963 4981
rect 44174 4972 44180 5024
rect 44232 5012 44238 5024
rect 44913 5015 44971 5021
rect 44913 5012 44925 5015
rect 44232 4984 44925 5012
rect 44232 4972 44238 4984
rect 44913 4981 44925 4984
rect 44959 4981 44971 5015
rect 44913 4975 44971 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 44542 4808 44548 4820
rect 44503 4780 44548 4808
rect 44542 4768 44548 4780
rect 44600 4768 44606 4820
rect 48130 4740 48136 4752
rect 44468 4712 48136 4740
rect 2958 4672 2964 4684
rect 2919 4644 2964 4672
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4295 4576 4721 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 7064 4576 7205 4604
rect 7064 4564 7070 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 40034 4564 40040 4616
rect 40092 4604 40098 4616
rect 40221 4607 40279 4613
rect 40221 4604 40233 4607
rect 40092 4576 40233 4604
rect 40092 4564 40098 4576
rect 40221 4573 40233 4576
rect 40267 4573 40279 4607
rect 40221 4567 40279 4573
rect 44266 4564 44272 4616
rect 44324 4604 44330 4616
rect 44468 4613 44496 4712
rect 48130 4700 48136 4712
rect 48188 4700 48194 4752
rect 46477 4675 46535 4681
rect 46477 4641 46489 4675
rect 46523 4672 46535 4675
rect 47946 4672 47952 4684
rect 46523 4644 47952 4672
rect 46523 4641 46535 4644
rect 46477 4635 46535 4641
rect 47946 4632 47952 4644
rect 48004 4632 48010 4684
rect 44453 4607 44511 4613
rect 44453 4604 44465 4607
rect 44324 4576 44465 4604
rect 44324 4564 44330 4576
rect 44453 4573 44465 4576
rect 44499 4573 44511 4607
rect 45186 4604 45192 4616
rect 45147 4576 45192 4604
rect 44453 4567 44511 4573
rect 45186 4564 45192 4576
rect 45244 4564 45250 4616
rect 45738 4564 45744 4616
rect 45796 4604 45802 4616
rect 45833 4607 45891 4613
rect 45833 4604 45845 4607
rect 45796 4576 45845 4604
rect 45796 4564 45802 4576
rect 45833 4573 45845 4576
rect 45879 4573 45891 4607
rect 45833 4567 45891 4573
rect 1762 4536 1768 4548
rect 1723 4508 1768 4536
rect 1762 4496 1768 4508
rect 1820 4496 1826 4548
rect 46474 4496 46480 4548
rect 46532 4536 46538 4548
rect 46661 4539 46719 4545
rect 46661 4536 46673 4539
rect 46532 4508 46673 4536
rect 46532 4496 46538 4508
rect 46661 4505 46673 4508
rect 46707 4505 46719 4539
rect 48314 4536 48320 4548
rect 48275 4508 48320 4536
rect 46661 4499 46719 4505
rect 48314 4496 48320 4508
rect 48372 4496 48378 4548
rect 45281 4471 45339 4477
rect 45281 4437 45293 4471
rect 45327 4468 45339 4471
rect 45370 4468 45376 4480
rect 45327 4440 45376 4468
rect 45327 4437 45339 4440
rect 45281 4431 45339 4437
rect 45370 4428 45376 4440
rect 45428 4428 45434 4480
rect 45830 4428 45836 4480
rect 45888 4468 45894 4480
rect 45925 4471 45983 4477
rect 45925 4468 45937 4471
rect 45888 4440 45937 4468
rect 45888 4428 45894 4440
rect 45925 4437 45937 4440
rect 45971 4437 45983 4471
rect 45925 4431 45983 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 2593 4267 2651 4273
rect 2593 4264 2605 4267
rect 1820 4236 2605 4264
rect 1820 4224 1826 4236
rect 2593 4233 2605 4236
rect 2639 4233 2651 4267
rect 2593 4227 2651 4233
rect 3804 4168 5212 4196
rect 1578 4088 1584 4140
rect 1636 4128 1642 4140
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1636 4100 2053 4128
rect 1636 4088 1642 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4097 2559 4131
rect 3142 4128 3148 4140
rect 3103 4100 3148 4128
rect 2501 4091 2559 4097
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 2516 4060 2544 4091
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3804 4128 3832 4168
rect 3712 4100 3832 4128
rect 5184 4128 5212 4168
rect 10244 4168 10548 4196
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 5184 4100 7021 4128
rect 3712 4060 3740 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 8294 4128 8300 4140
rect 8207 4100 8300 4128
rect 7009 4091 7067 4097
rect 2004 4032 3740 4060
rect 2004 4020 2010 4032
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 3844 4032 3889 4060
rect 3844 4020 3850 4032
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 4249 4063 4307 4069
rect 4028 4032 4073 4060
rect 4028 4020 4034 4032
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 7024 4060 7052 4091
rect 8294 4088 8300 4100
rect 8352 4128 8358 4140
rect 10244 4128 10272 4168
rect 10410 4128 10416 4140
rect 8352 4100 10272 4128
rect 10371 4100 10416 4128
rect 8352 4088 8358 4100
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 10520 4128 10548 4168
rect 38672 4168 40080 4196
rect 10520 4100 12434 4128
rect 10594 4060 10600 4072
rect 7024 4032 10600 4060
rect 4249 4023 4307 4029
rect 4062 3952 4068 4004
rect 4120 3992 4126 4004
rect 4264 3992 4292 4023
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 12406 4060 12434 4100
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12952 4100 13001 4128
rect 12952 4088 12958 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 38672 4128 38700 4168
rect 12989 4091 13047 4097
rect 26206 4100 38700 4128
rect 40052 4128 40080 4168
rect 43717 4131 43775 4137
rect 43717 4128 43729 4131
rect 40052 4100 43729 4128
rect 20714 4060 20720 4072
rect 12406 4032 20720 4060
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 4120 3964 4292 3992
rect 4120 3952 4126 3964
rect 12894 3952 12900 4004
rect 12952 3992 12958 4004
rect 26206 3992 26234 4100
rect 43717 4097 43729 4100
rect 43763 4097 43775 4131
rect 44358 4128 44364 4140
rect 44319 4100 44364 4128
rect 43717 4091 43775 4097
rect 38654 4060 38660 4072
rect 38615 4032 38660 4060
rect 38654 4020 38660 4032
rect 38712 4020 38718 4072
rect 38841 4063 38899 4069
rect 38841 4029 38853 4063
rect 38887 4060 38899 4063
rect 39390 4060 39396 4072
rect 38887 4032 39396 4060
rect 38887 4029 38899 4032
rect 38841 4023 38899 4029
rect 39390 4020 39396 4032
rect 39448 4020 39454 4072
rect 39485 4063 39543 4069
rect 39485 4029 39497 4063
rect 39531 4029 39543 4063
rect 39485 4023 39543 4029
rect 12952 3964 26234 3992
rect 12952 3952 12958 3964
rect 39298 3952 39304 4004
rect 39356 3992 39362 4004
rect 39500 3992 39528 4023
rect 39356 3964 39528 3992
rect 43732 3992 43760 4091
rect 44358 4088 44364 4100
rect 44416 4088 44422 4140
rect 47946 4128 47952 4140
rect 47907 4100 47952 4128
rect 47946 4088 47952 4100
rect 48004 4088 48010 4140
rect 45373 4063 45431 4069
rect 45373 4029 45385 4063
rect 45419 4029 45431 4063
rect 45373 4023 45431 4029
rect 45557 4063 45615 4069
rect 45557 4029 45569 4063
rect 45603 4060 45615 4063
rect 46934 4060 46940 4072
rect 45603 4032 46940 4060
rect 45603 4029 45615 4032
rect 45557 4023 45615 4029
rect 45388 3992 45416 4023
rect 46934 4020 46940 4032
rect 46992 4020 46998 4072
rect 47213 4063 47271 4069
rect 47213 4029 47225 4063
rect 47259 4060 47271 4063
rect 47670 4060 47676 4072
rect 47259 4032 47676 4060
rect 47259 4029 47271 4032
rect 47213 4023 47271 4029
rect 47670 4020 47676 4032
rect 47728 4020 47734 4072
rect 47946 3992 47952 4004
rect 43732 3964 45232 3992
rect 45388 3964 47952 3992
rect 39356 3952 39362 3964
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3970 3924 3976 3936
rect 3283 3896 3976 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7101 3927 7159 3933
rect 7101 3924 7113 3927
rect 6972 3896 7113 3924
rect 6972 3884 6978 3896
rect 7101 3893 7113 3896
rect 7147 3893 7159 3927
rect 7101 3887 7159 3893
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7616 3896 7849 3924
rect 7616 3884 7622 3896
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 8386 3924 8392 3936
rect 8347 3896 8392 3924
rect 7837 3887 7895 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12526 3924 12532 3936
rect 12483 3896 12532 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 13081 3927 13139 3933
rect 13081 3893 13093 3927
rect 13127 3924 13139 3927
rect 13170 3924 13176 3936
rect 13127 3896 13176 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 24762 3884 24768 3936
rect 24820 3924 24826 3936
rect 25409 3927 25467 3933
rect 25409 3924 25421 3927
rect 24820 3896 25421 3924
rect 24820 3884 24826 3896
rect 25409 3893 25421 3896
rect 25455 3893 25467 3927
rect 25409 3887 25467 3893
rect 25866 3884 25872 3936
rect 25924 3924 25930 3936
rect 26145 3927 26203 3933
rect 26145 3924 26157 3927
rect 25924 3896 26157 3924
rect 25924 3884 25930 3896
rect 26145 3893 26157 3896
rect 26191 3893 26203 3927
rect 26145 3887 26203 3893
rect 40494 3884 40500 3936
rect 40552 3924 40558 3936
rect 41141 3927 41199 3933
rect 41141 3924 41153 3927
rect 40552 3896 41153 3924
rect 40552 3884 40558 3896
rect 41141 3893 41153 3896
rect 41187 3893 41199 3927
rect 41141 3887 41199 3893
rect 41785 3927 41843 3933
rect 41785 3893 41797 3927
rect 41831 3924 41843 3927
rect 42610 3924 42616 3936
rect 41831 3896 42616 3924
rect 41831 3893 41843 3896
rect 41785 3887 41843 3893
rect 42610 3884 42616 3896
rect 42668 3884 42674 3936
rect 42978 3884 42984 3936
rect 43036 3924 43042 3936
rect 43809 3927 43867 3933
rect 43809 3924 43821 3927
rect 43036 3896 43821 3924
rect 43036 3884 43042 3896
rect 43809 3893 43821 3896
rect 43855 3893 43867 3927
rect 43809 3887 43867 3893
rect 44453 3927 44511 3933
rect 44453 3893 44465 3927
rect 44499 3924 44511 3927
rect 45094 3924 45100 3936
rect 44499 3896 45100 3924
rect 44499 3893 44511 3896
rect 44453 3887 44511 3893
rect 45094 3884 45100 3896
rect 45152 3884 45158 3936
rect 45204 3924 45232 3964
rect 47946 3952 47952 3964
rect 48004 3952 48010 4004
rect 47762 3924 47768 3936
rect 45204 3896 47768 3924
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 4706 3720 4712 3732
rect 1688 3692 4712 3720
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1688 3584 1716 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 5534 3720 5540 3732
rect 4856 3692 5540 3720
rect 4856 3680 4862 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6012 3692 6224 3720
rect 5350 3652 5356 3664
rect 1780 3624 5356 3652
rect 1780 3593 1808 3624
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 6012 3652 6040 3692
rect 5552 3624 6040 3652
rect 5552 3600 5580 3624
rect 1627 3556 1716 3584
rect 1765 3587 1823 3593
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1765 3553 1777 3587
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 2832 3556 2877 3584
rect 2832 3544 2838 3556
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3970 3584 3976 3596
rect 3200 3556 3976 3584
rect 3200 3544 3206 3556
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3584 5135 3587
rect 5460 3584 5580 3600
rect 6196 3593 6224 3692
rect 24578 3680 24584 3732
rect 24636 3720 24642 3732
rect 44358 3720 44364 3732
rect 24636 3692 44364 3720
rect 24636 3680 24642 3692
rect 44358 3680 44364 3692
rect 44416 3680 44422 3732
rect 47026 3652 47032 3664
rect 12406 3624 19472 3652
rect 5123 3572 5580 3584
rect 6181 3587 6239 3593
rect 5123 3556 5488 3572
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 6181 3553 6193 3587
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6512 3556 6653 3584
rect 6512 3544 6518 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 10502 3584 10508 3596
rect 10463 3556 10508 3584
rect 6641 3547 6699 3553
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4212 3488 4445 3516
rect 4212 3476 4218 3488
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 10318 3516 10324 3528
rect 10279 3488 10324 3516
rect 5537 3479 5595 3485
rect 2590 3408 2596 3460
rect 2648 3448 2654 3460
rect 5552 3448 5580 3479
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 2648 3420 5580 3448
rect 2648 3408 2654 3420
rect 5552 3380 5580 3420
rect 5629 3451 5687 3457
rect 5629 3417 5641 3451
rect 5675 3448 5687 3451
rect 6365 3451 6423 3457
rect 6365 3448 6377 3451
rect 5675 3420 6377 3448
rect 5675 3417 5687 3420
rect 5629 3411 5687 3417
rect 6365 3417 6377 3420
rect 6411 3417 6423 3451
rect 6365 3411 6423 3417
rect 12406 3380 12434 3624
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13173 3519 13231 3525
rect 13173 3516 13185 3519
rect 13044 3488 13185 3516
rect 13044 3476 13050 3488
rect 13173 3485 13185 3488
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16908 3488 16957 3516
rect 16908 3476 16914 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 17402 3516 17408 3528
rect 17315 3488 17408 3516
rect 16945 3479 17003 3485
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 19334 3516 19340 3528
rect 18923 3488 19340 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19444 3525 19472 3624
rect 25148 3624 47032 3652
rect 25148 3584 25176 3624
rect 47026 3612 47032 3624
rect 47084 3612 47090 3664
rect 25866 3584 25872 3596
rect 20732 3556 25176 3584
rect 25827 3556 25872 3584
rect 20732 3528 20760 3556
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 20254 3516 20260 3528
rect 20215 3488 20260 3516
rect 19429 3479 19487 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20714 3516 20720 3528
rect 20675 3488 20720 3516
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 22002 3476 22008 3528
rect 22060 3516 22066 3528
rect 22664 3525 22692 3556
rect 25866 3544 25872 3556
rect 25924 3544 25930 3596
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 39390 3584 39396 3596
rect 39351 3556 39396 3584
rect 39390 3544 39396 3556
rect 39448 3544 39454 3596
rect 40494 3584 40500 3596
rect 40455 3556 40500 3584
rect 40494 3544 40500 3556
rect 40552 3544 40558 3596
rect 41230 3584 41236 3596
rect 41191 3556 41236 3584
rect 41230 3544 41236 3556
rect 41288 3544 41294 3596
rect 44266 3584 44272 3596
rect 42812 3556 44272 3584
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 22060 3488 22201 3516
rect 22060 3476 22066 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 22649 3519 22707 3525
rect 22649 3485 22661 3519
rect 22695 3485 22707 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 22649 3479 22707 3485
rect 24578 3476 24584 3488
rect 24636 3516 24642 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 24636 3488 25237 3516
rect 24636 3476 24642 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 27430 3476 27436 3528
rect 27488 3516 27494 3528
rect 28353 3519 28411 3525
rect 28353 3516 28365 3519
rect 27488 3488 28365 3516
rect 27488 3476 27494 3488
rect 28353 3485 28365 3488
rect 28399 3485 28411 3519
rect 31846 3516 31852 3528
rect 31807 3488 31852 3516
rect 28353 3479 28411 3485
rect 31846 3476 31852 3488
rect 31904 3476 31910 3528
rect 32306 3516 32312 3528
rect 32219 3488 32312 3516
rect 32306 3476 32312 3488
rect 32364 3516 32370 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 32364 3488 38025 3516
rect 32364 3476 32370 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 38841 3519 38899 3525
rect 38841 3516 38853 3519
rect 38436 3488 38853 3516
rect 38436 3476 38442 3488
rect 38841 3485 38853 3488
rect 38887 3485 38899 3519
rect 38841 3479 38899 3485
rect 39301 3519 39359 3525
rect 39301 3485 39313 3519
rect 39347 3485 39359 3519
rect 39301 3479 39359 3485
rect 17420 3448 17448 3476
rect 25317 3451 25375 3457
rect 17420 3420 25084 3448
rect 5552 3352 12434 3380
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 17092 3352 17509 3380
rect 17092 3340 17098 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 17497 3343 17555 3349
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 19484 3352 19533 3380
rect 19484 3340 19490 3352
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 20806 3380 20812 3392
rect 20767 3352 20812 3380
rect 19521 3343 19579 3349
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 22186 3340 22192 3392
rect 22244 3380 22250 3392
rect 22741 3383 22799 3389
rect 22741 3380 22753 3383
rect 22244 3352 22753 3380
rect 22244 3340 22250 3352
rect 22741 3349 22753 3352
rect 22787 3349 22799 3383
rect 22741 3343 22799 3349
rect 24673 3383 24731 3389
rect 24673 3349 24685 3383
rect 24719 3380 24731 3383
rect 24946 3380 24952 3392
rect 24719 3352 24952 3380
rect 24719 3349 24731 3352
rect 24673 3343 24731 3349
rect 24946 3340 24952 3352
rect 25004 3340 25010 3392
rect 25056 3380 25084 3420
rect 25317 3417 25329 3451
rect 25363 3448 25375 3451
rect 26053 3451 26111 3457
rect 26053 3448 26065 3451
rect 25363 3420 26065 3448
rect 25363 3417 25375 3420
rect 25317 3411 25375 3417
rect 26053 3417 26065 3420
rect 26099 3417 26111 3451
rect 26053 3411 26111 3417
rect 27522 3380 27528 3392
rect 25056 3352 27528 3380
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 32401 3383 32459 3389
rect 32401 3349 32413 3383
rect 32447 3380 32459 3383
rect 32490 3380 32496 3392
rect 32447 3352 32496 3380
rect 32447 3349 32459 3352
rect 32401 3343 32459 3349
rect 32490 3340 32496 3352
rect 32548 3340 32554 3392
rect 38105 3383 38163 3389
rect 38105 3349 38117 3383
rect 38151 3380 38163 3383
rect 38562 3380 38568 3392
rect 38151 3352 38568 3380
rect 38151 3349 38163 3352
rect 38105 3343 38163 3349
rect 38562 3340 38568 3352
rect 38620 3340 38626 3392
rect 39316 3380 39344 3479
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 42812 3525 42840 3556
rect 44266 3544 44272 3556
rect 44324 3544 44330 3596
rect 45649 3587 45707 3593
rect 45649 3553 45661 3587
rect 45695 3584 45707 3587
rect 48133 3587 48191 3593
rect 48133 3584 48145 3587
rect 45695 3556 48145 3584
rect 45695 3553 45707 3556
rect 45649 3547 45707 3553
rect 48133 3553 48145 3556
rect 48179 3553 48191 3587
rect 48133 3547 48191 3553
rect 42797 3519 42855 3525
rect 42797 3516 42809 3519
rect 42484 3488 42809 3516
rect 42484 3476 42490 3488
rect 42797 3485 42809 3488
rect 42843 3485 42855 3519
rect 42797 3479 42855 3485
rect 43901 3519 43959 3525
rect 43901 3485 43913 3519
rect 43947 3516 43959 3519
rect 44450 3516 44456 3528
rect 43947 3488 44456 3516
rect 43947 3485 43959 3488
rect 43901 3479 43959 3485
rect 44450 3476 44456 3488
rect 44508 3476 44514 3528
rect 44545 3519 44603 3525
rect 44545 3485 44557 3519
rect 44591 3516 44603 3519
rect 44910 3516 44916 3528
rect 44591 3488 44916 3516
rect 44591 3485 44603 3488
rect 44545 3479 44603 3485
rect 44910 3476 44916 3488
rect 44968 3476 44974 3528
rect 40681 3451 40739 3457
rect 40681 3417 40693 3451
rect 40727 3448 40739 3451
rect 41414 3448 41420 3460
rect 40727 3420 41420 3448
rect 40727 3417 40739 3420
rect 40681 3411 40739 3417
rect 41414 3408 41420 3420
rect 41472 3408 41478 3460
rect 45830 3448 45836 3460
rect 42444 3420 45554 3448
rect 45791 3420 45836 3448
rect 42444 3380 42472 3420
rect 39316 3352 42472 3380
rect 42794 3340 42800 3392
rect 42852 3380 42858 3392
rect 42889 3383 42947 3389
rect 42889 3380 42901 3383
rect 42852 3352 42901 3380
rect 42852 3340 42858 3352
rect 42889 3349 42901 3352
rect 42935 3349 42947 3383
rect 45526 3380 45554 3420
rect 45830 3408 45836 3420
rect 45888 3408 45894 3460
rect 47026 3408 47032 3460
rect 47084 3448 47090 3460
rect 47489 3451 47547 3457
rect 47489 3448 47501 3451
rect 47084 3420 47501 3448
rect 47084 3408 47090 3420
rect 47489 3417 47501 3420
rect 47535 3417 47547 3451
rect 47489 3411 47547 3417
rect 47394 3380 47400 3392
rect 45526 3352 47400 3380
rect 42889 3343 42947 3349
rect 47394 3340 47400 3352
rect 47452 3340 47458 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 4982 3176 4988 3188
rect 2746 3148 4988 3176
rect 2746 3108 2774 3148
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 45738 3176 45744 3188
rect 40696 3148 45744 3176
rect 1872 3080 2774 3108
rect 4341 3111 4399 3117
rect 1872 3049 1900 3080
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 5626 3108 5632 3120
rect 4387 3080 5632 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 7745 3111 7803 3117
rect 7745 3077 7757 3111
rect 7791 3108 7803 3111
rect 8386 3108 8392 3120
rect 7791 3080 8392 3108
rect 7791 3077 7803 3080
rect 7745 3071 7803 3077
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 13170 3108 13176 3120
rect 13131 3080 13176 3108
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 17034 3108 17040 3120
rect 16995 3080 17040 3108
rect 17034 3068 17040 3080
rect 17092 3068 17098 3120
rect 19797 3111 19855 3117
rect 19797 3077 19809 3111
rect 19843 3108 19855 3111
rect 20806 3108 20812 3120
rect 19843 3080 20812 3108
rect 19843 3077 19855 3080
rect 19797 3071 19855 3077
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 22186 3108 22192 3120
rect 22147 3080 22192 3108
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 24946 3108 24952 3120
rect 24907 3080 24952 3108
rect 24946 3068 24952 3080
rect 25004 3068 25010 3120
rect 32490 3108 32496 3120
rect 32451 3080 32496 3108
rect 32490 3068 32496 3080
rect 32548 3068 32554 3120
rect 38562 3108 38568 3120
rect 38523 3080 38568 3108
rect 38562 3068 38568 3080
rect 38620 3068 38626 3120
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 1857 3003 1915 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 7558 3040 7564 3052
rect 7519 3012 7564 3040
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 10376 3012 10517 3040
rect 10376 3000 10382 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 10652 3012 12357 3040
rect 10652 3000 10658 3012
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12345 3003 12403 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 24762 3040 24768 3052
rect 24723 3012 24768 3040
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 27430 3040 27436 3052
rect 27391 3012 27436 3040
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 31846 3000 31852 3052
rect 31904 3040 31910 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31904 3012 32321 3040
rect 31904 3000 31910 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 38378 3040 38384 3052
rect 38339 3012 38384 3040
rect 32309 3003 32367 3009
rect 38378 3000 38384 3012
rect 38436 3000 38442 3052
rect 40696 3049 40724 3148
rect 45738 3136 45744 3148
rect 45796 3136 45802 3188
rect 41414 3108 41420 3120
rect 41375 3080 41420 3108
rect 41414 3068 41420 3080
rect 41472 3068 41478 3120
rect 42794 3108 42800 3120
rect 42755 3080 42800 3108
rect 42794 3068 42800 3080
rect 42852 3068 42858 3120
rect 45094 3108 45100 3120
rect 45055 3080 45100 3108
rect 45094 3068 45100 3080
rect 45152 3068 45158 3120
rect 40681 3043 40739 3049
rect 40681 3009 40693 3043
rect 40727 3009 40739 3043
rect 40681 3003 40739 3009
rect 41325 3043 41383 3049
rect 41325 3009 41337 3043
rect 41371 3040 41383 3043
rect 42426 3040 42432 3052
rect 41371 3012 42432 3040
rect 41371 3009 41383 3012
rect 41325 3003 41383 3009
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 42610 3040 42616 3052
rect 42571 3012 42616 3040
rect 42610 3000 42616 3012
rect 42668 3000 42674 3052
rect 44910 3040 44916 3052
rect 44871 3012 44916 3040
rect 44910 3000 44916 3012
rect 44968 3000 44974 3052
rect 47946 3040 47952 3052
rect 47907 3012 47952 3040
rect 47946 3000 47952 3012
rect 48004 3000 48010 3052
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2941 2099 2975
rect 2866 2972 2872 2984
rect 2827 2944 2872 2972
rect 2041 2935 2099 2941
rect 2056 2904 2084 2935
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7892 2944 8033 2972
rect 7892 2932 7898 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 13538 2972 13544 2984
rect 13499 2944 13544 2972
rect 8021 2935 8079 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 17402 2972 17408 2984
rect 17363 2944 17408 2972
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2972 19671 2975
rect 20254 2972 20260 2984
rect 19659 2944 20260 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 25774 2972 25780 2984
rect 25735 2944 25780 2972
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 27614 2972 27620 2984
rect 27575 2944 27620 2972
rect 27614 2932 27620 2944
rect 27672 2932 27678 2984
rect 27706 2932 27712 2984
rect 27764 2972 27770 2984
rect 27893 2975 27951 2981
rect 27893 2972 27905 2975
rect 27764 2944 27905 2972
rect 27764 2932 27770 2944
rect 27893 2941 27905 2944
rect 27939 2941 27951 2975
rect 27893 2935 27951 2941
rect 32214 2932 32220 2984
rect 32272 2972 32278 2984
rect 32769 2975 32827 2981
rect 32769 2972 32781 2975
rect 32272 2944 32781 2972
rect 32272 2932 32278 2944
rect 32769 2941 32781 2944
rect 32815 2941 32827 2975
rect 32769 2935 32827 2941
rect 40221 2975 40279 2981
rect 40221 2941 40233 2975
rect 40267 2941 40279 2975
rect 40221 2935 40279 2941
rect 4706 2904 4712 2916
rect 2056 2876 4712 2904
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 40236 2904 40264 2935
rect 41874 2932 41880 2984
rect 41932 2972 41938 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 41932 2944 43085 2972
rect 41932 2932 41938 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 45094 2932 45100 2984
rect 45152 2972 45158 2984
rect 45373 2975 45431 2981
rect 45373 2972 45385 2975
rect 45152 2944 45385 2972
rect 45152 2932 45158 2944
rect 45373 2941 45385 2944
rect 45419 2941 45431 2975
rect 45373 2935 45431 2941
rect 46750 2904 46756 2916
rect 40236 2876 46756 2904
rect 46750 2864 46756 2876
rect 46808 2864 46814 2916
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 4062 2836 4068 2848
rect 3292 2808 4068 2836
rect 3292 2796 3298 2808
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 7098 2836 7104 2848
rect 7059 2808 7104 2836
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 12434 2836 12440 2848
rect 12395 2808 12440 2836
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 40218 2796 40224 2848
rect 40276 2836 40282 2848
rect 40773 2839 40831 2845
rect 40773 2836 40785 2839
rect 40276 2808 40785 2836
rect 40276 2796 40282 2808
rect 40773 2805 40785 2808
rect 40819 2805 40831 2839
rect 40773 2799 40831 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 4157 2635 4215 2641
rect 4157 2632 4169 2635
rect 3844 2604 4169 2632
rect 3844 2592 3850 2604
rect 4157 2601 4169 2604
rect 4203 2601 4215 2635
rect 4157 2595 4215 2601
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5626 2632 5632 2644
rect 4764 2604 4809 2632
rect 5587 2604 5632 2632
rect 4764 2592 4770 2604
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 12894 2632 12900 2644
rect 6886 2604 12900 2632
rect 5718 2524 5724 2576
rect 5776 2564 5782 2576
rect 6886 2564 6914 2604
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 27614 2632 27620 2644
rect 27575 2604 27620 2632
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 38654 2592 38660 2644
rect 38712 2632 38718 2644
rect 38933 2635 38991 2641
rect 38933 2632 38945 2635
rect 38712 2604 38945 2632
rect 38712 2592 38718 2604
rect 38933 2601 38945 2604
rect 38979 2601 38991 2635
rect 38933 2595 38991 2601
rect 46934 2592 46940 2644
rect 46992 2632 46998 2644
rect 47857 2635 47915 2641
rect 47857 2632 47869 2635
rect 46992 2604 47869 2632
rect 46992 2592 46998 2604
rect 47857 2601 47869 2604
rect 47903 2601 47915 2635
rect 47857 2595 47915 2601
rect 12526 2564 12532 2576
rect 5776 2536 6914 2564
rect 11900 2536 12532 2564
rect 5776 2524 5782 2536
rect 658 2456 664 2508
rect 716 2496 722 2508
rect 2041 2499 2099 2505
rect 2041 2496 2053 2499
rect 716 2468 2053 2496
rect 716 2456 722 2468
rect 2041 2465 2053 2468
rect 2087 2465 2099 2499
rect 2041 2459 2099 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7098 2496 7104 2508
rect 6779 2468 7104 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 11900 2505 11928 2536
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 19426 2524 19432 2576
rect 19484 2524 19490 2576
rect 44174 2564 44180 2576
rect 42812 2536 44180 2564
rect 11885 2499 11943 2505
rect 7248 2468 7293 2496
rect 7248 2456 7254 2468
rect 11885 2465 11897 2499
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 12069 2499 12127 2505
rect 12069 2465 12081 2499
rect 12115 2496 12127 2499
rect 12434 2496 12440 2508
rect 12115 2468 12440 2496
rect 12115 2465 12127 2468
rect 12069 2459 12127 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 12894 2496 12900 2508
rect 12855 2468 12900 2496
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 19444 2496 19472 2524
rect 19613 2499 19671 2505
rect 19613 2496 19625 2499
rect 19444 2468 19625 2496
rect 19613 2465 19625 2468
rect 19659 2465 19671 2499
rect 19613 2459 19671 2465
rect 19702 2456 19708 2508
rect 19760 2496 19766 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19760 2468 19901 2496
rect 19760 2456 19766 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 24302 2456 24308 2508
rect 24360 2496 24366 2508
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 24360 2468 24869 2496
rect 24360 2456 24366 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 40034 2496 40040 2508
rect 39995 2468 40040 2496
rect 24857 2459 24915 2465
rect 40034 2456 40040 2468
rect 40092 2456 40098 2508
rect 40218 2496 40224 2508
rect 40179 2468 40224 2496
rect 40218 2456 40224 2468
rect 40276 2456 40282 2508
rect 40586 2496 40592 2508
rect 40547 2468 40592 2496
rect 40586 2456 40592 2468
rect 40644 2456 40650 2508
rect 42812 2505 42840 2536
rect 44174 2524 44180 2536
rect 44232 2524 44238 2576
rect 42797 2499 42855 2505
rect 42797 2465 42809 2499
rect 42843 2465 42855 2499
rect 42978 2496 42984 2508
rect 42939 2468 42984 2496
rect 42797 2459 42855 2465
rect 42978 2456 42984 2468
rect 43036 2456 43042 2508
rect 44450 2456 44456 2508
rect 44508 2496 44514 2508
rect 45189 2499 45247 2505
rect 45189 2496 45201 2499
rect 44508 2468 45201 2496
rect 44508 2456 44514 2468
rect 45189 2465 45201 2468
rect 45235 2465 45247 2499
rect 45370 2496 45376 2508
rect 45331 2468 45376 2496
rect 45189 2459 45247 2465
rect 45370 2456 45376 2468
rect 45428 2456 45434 2508
rect 45738 2496 45744 2508
rect 45699 2468 45744 2496
rect 45738 2456 45744 2468
rect 45796 2456 45802 2508
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1596 2292 1624 2391
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4212 2400 4629 2428
rect 4212 2388 4218 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2428 5595 2431
rect 5718 2428 5724 2440
rect 5583 2400 5724 2428
rect 5583 2397 5595 2400
rect 5537 2391 5595 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19392 2400 19441 2428
rect 19392 2388 19398 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23900 2400 24593 2428
rect 23900 2388 23906 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 27522 2428 27528 2440
rect 27435 2400 27528 2428
rect 24581 2391 24639 2397
rect 27522 2388 27528 2400
rect 27580 2428 27586 2440
rect 32306 2428 32312 2440
rect 27580 2400 32312 2428
rect 27580 2388 27586 2400
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 47762 2428 47768 2440
rect 47723 2400 47768 2428
rect 47762 2388 47768 2400
rect 47820 2388 47826 2440
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2360 1823 2363
rect 4890 2360 4896 2372
rect 1811 2332 4896 2360
rect 1811 2329 1823 2332
rect 1765 2323 1823 2329
rect 4890 2320 4896 2332
rect 4948 2320 4954 2372
rect 6914 2320 6920 2372
rect 6972 2360 6978 2372
rect 44637 2363 44695 2369
rect 6972 2332 7017 2360
rect 6972 2320 6978 2332
rect 44637 2329 44649 2363
rect 44683 2329 44695 2363
rect 44637 2323 44695 2329
rect 7006 2292 7012 2304
rect 1596 2264 7012 2292
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 44652 2292 44680 2323
rect 46842 2292 46848 2304
rect 44652 2264 46848 2292
rect 46842 2252 46848 2264
rect 46900 2252 46906 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
<< via1 >>
rect 20 48764 72 48816
rect 8024 48764 8076 48816
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 4896 47132 4948 47184
rect 3516 47064 3568 47116
rect 7012 47064 7064 47116
rect 47216 47107 47268 47116
rect 47216 47073 47225 47107
rect 47225 47073 47259 47107
rect 47259 47073 47268 47107
rect 47216 47064 47268 47073
rect 2044 46996 2096 47048
rect 2688 47039 2740 47048
rect 2688 47005 2697 47039
rect 2697 47005 2731 47039
rect 2731 47005 2740 47039
rect 2688 46996 2740 47005
rect 4160 46996 4212 47048
rect 5540 46996 5592 47048
rect 5724 46996 5776 47048
rect 6552 46996 6604 47048
rect 7380 47039 7432 47048
rect 7380 47005 7389 47039
rect 7389 47005 7423 47039
rect 7423 47005 7432 47039
rect 7380 46996 7432 47005
rect 8024 47039 8076 47048
rect 8024 47005 8033 47039
rect 8033 47005 8067 47039
rect 8067 47005 8076 47039
rect 8024 46996 8076 47005
rect 8392 46996 8444 47048
rect 12532 47039 12584 47048
rect 12532 47005 12541 47039
rect 12541 47005 12575 47039
rect 12575 47005 12584 47039
rect 12532 46996 12584 47005
rect 14556 47039 14608 47048
rect 14556 47005 14565 47039
rect 14565 47005 14599 47039
rect 14599 47005 14608 47039
rect 14556 46996 14608 47005
rect 15200 47039 15252 47048
rect 15200 47005 15209 47039
rect 15209 47005 15243 47039
rect 15243 47005 15252 47039
rect 15200 46996 15252 47005
rect 22468 46996 22520 47048
rect 25320 47039 25372 47048
rect 25320 47005 25329 47039
rect 25329 47005 25363 47039
rect 25363 47005 25372 47039
rect 25320 46996 25372 47005
rect 27160 46996 27212 47048
rect 27988 47039 28040 47048
rect 27988 47005 27997 47039
rect 27997 47005 28031 47039
rect 28031 47005 28040 47039
rect 27988 46996 28040 47005
rect 29092 47039 29144 47048
rect 29092 47005 29101 47039
rect 29101 47005 29135 47039
rect 29135 47005 29144 47039
rect 29092 46996 29144 47005
rect 29920 47039 29972 47048
rect 29920 47005 29929 47039
rect 29929 47005 29963 47039
rect 29963 47005 29972 47039
rect 29920 46996 29972 47005
rect 33232 47039 33284 47048
rect 33232 47005 33241 47039
rect 33241 47005 33275 47039
rect 33275 47005 33284 47039
rect 33232 46996 33284 47005
rect 39764 46996 39816 47048
rect 42616 46996 42668 47048
rect 44640 47039 44692 47048
rect 44640 47005 44649 47039
rect 44649 47005 44683 47039
rect 44683 47005 44692 47039
rect 44640 46996 44692 47005
rect 45376 47039 45428 47048
rect 45376 47005 45385 47039
rect 45385 47005 45419 47039
rect 45419 47005 45428 47039
rect 45376 46996 45428 47005
rect 47676 46996 47728 47048
rect 4804 46928 4856 46980
rect 45560 46971 45612 46980
rect 45560 46937 45569 46971
rect 45569 46937 45603 46971
rect 45603 46937 45612 46971
rect 47860 46971 47912 46980
rect 45560 46928 45612 46937
rect 47860 46937 47869 46971
rect 47869 46937 47903 46971
rect 47903 46937 47912 46971
rect 47860 46928 47912 46937
rect 1768 46860 1820 46912
rect 6736 46860 6788 46912
rect 7840 46903 7892 46912
rect 7840 46869 7849 46903
rect 7849 46869 7883 46903
rect 7883 46869 7892 46903
rect 7840 46860 7892 46869
rect 9128 46903 9180 46912
rect 9128 46869 9137 46903
rect 9137 46869 9171 46903
rect 9171 46869 9180 46903
rect 9128 46860 9180 46869
rect 27804 46903 27856 46912
rect 27804 46869 27813 46903
rect 27813 46869 27847 46903
rect 27847 46869 27856 46903
rect 27804 46860 27856 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 7380 46656 7432 46708
rect 4068 46588 4120 46640
rect 6736 46631 6788 46640
rect 6736 46597 6745 46631
rect 6745 46597 6779 46631
rect 6779 46597 6788 46631
rect 6736 46588 6788 46597
rect 4160 46563 4212 46572
rect 4160 46529 4169 46563
rect 4169 46529 4203 46563
rect 4203 46529 4212 46563
rect 4160 46520 4212 46529
rect 6552 46563 6604 46572
rect 6552 46529 6561 46563
rect 6561 46529 6595 46563
rect 6595 46529 6604 46563
rect 6552 46520 6604 46529
rect 12532 46588 12584 46640
rect 15200 46588 15252 46640
rect 22468 46563 22520 46572
rect 22468 46529 22477 46563
rect 22477 46529 22511 46563
rect 22511 46529 22520 46563
rect 22468 46520 22520 46529
rect 25320 46588 25372 46640
rect 27160 46563 27212 46572
rect 27160 46529 27169 46563
rect 27169 46529 27203 46563
rect 27203 46529 27212 46563
rect 27160 46520 27212 46529
rect 29092 46520 29144 46572
rect 33232 46588 33284 46640
rect 48320 46588 48372 46640
rect 39764 46563 39816 46572
rect 39764 46529 39773 46563
rect 39773 46529 39807 46563
rect 39807 46529 39816 46563
rect 39764 46520 39816 46529
rect 42616 46563 42668 46572
rect 42616 46529 42625 46563
rect 42625 46529 42659 46563
rect 42659 46529 42668 46563
rect 42616 46520 42668 46529
rect 44640 46520 44692 46572
rect 2596 46452 2648 46504
rect 4620 46452 4672 46504
rect 4712 46495 4764 46504
rect 4712 46461 4721 46495
rect 4721 46461 4755 46495
rect 4755 46461 4764 46495
rect 7012 46495 7064 46504
rect 4712 46452 4764 46461
rect 7012 46461 7021 46495
rect 7021 46461 7055 46495
rect 7055 46461 7064 46495
rect 7012 46452 7064 46461
rect 12440 46452 12492 46504
rect 12900 46495 12952 46504
rect 12900 46461 12909 46495
rect 12909 46461 12943 46495
rect 12943 46461 12952 46495
rect 12900 46452 12952 46461
rect 14648 46495 14700 46504
rect 14648 46461 14657 46495
rect 14657 46461 14691 46495
rect 14691 46461 14700 46495
rect 14648 46452 14700 46461
rect 15476 46495 15528 46504
rect 15476 46461 15485 46495
rect 15485 46461 15519 46495
rect 15519 46461 15528 46495
rect 15476 46452 15528 46461
rect 22928 46452 22980 46504
rect 23204 46495 23256 46504
rect 23204 46461 23213 46495
rect 23213 46461 23247 46495
rect 23247 46461 23256 46495
rect 23204 46452 23256 46461
rect 24952 46495 25004 46504
rect 24952 46461 24961 46495
rect 24961 46461 24995 46495
rect 24995 46461 25004 46495
rect 24952 46452 25004 46461
rect 25780 46495 25832 46504
rect 25780 46461 25789 46495
rect 25789 46461 25823 46495
rect 25823 46461 25832 46495
rect 25780 46452 25832 46461
rect 26976 46452 27028 46504
rect 29644 46495 29696 46504
rect 1952 46384 2004 46436
rect 2964 46384 3016 46436
rect 27068 46384 27120 46436
rect 29644 46461 29653 46495
rect 29653 46461 29687 46495
rect 29687 46461 29696 46495
rect 29644 46452 29696 46461
rect 29736 46452 29788 46504
rect 33232 46452 33284 46504
rect 33508 46495 33560 46504
rect 33508 46461 33517 46495
rect 33517 46461 33551 46495
rect 33551 46461 33560 46495
rect 33508 46452 33560 46461
rect 37648 46495 37700 46504
rect 37648 46461 37657 46495
rect 37657 46461 37691 46495
rect 37691 46461 37700 46495
rect 37648 46452 37700 46461
rect 39948 46495 40000 46504
rect 36728 46384 36780 46436
rect 39948 46461 39957 46495
rect 39957 46461 39991 46495
rect 39991 46461 40000 46495
rect 39948 46452 40000 46461
rect 42800 46495 42852 46504
rect 38660 46384 38712 46436
rect 42800 46461 42809 46495
rect 42809 46461 42843 46495
rect 42843 46461 42852 46495
rect 42800 46452 42852 46461
rect 41880 46384 41932 46436
rect 48044 46452 48096 46504
rect 10416 46316 10468 46368
rect 22744 46316 22796 46368
rect 29736 46316 29788 46368
rect 35532 46316 35584 46368
rect 45744 46316 45796 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 4896 46112 4948 46164
rect 22744 46112 22796 46164
rect 22928 46155 22980 46164
rect 22928 46121 22937 46155
rect 22937 46121 22971 46155
rect 22971 46121 22980 46155
rect 22928 46112 22980 46121
rect 26976 46155 27028 46164
rect 26976 46121 26985 46155
rect 26985 46121 27019 46155
rect 27019 46121 27028 46155
rect 26976 46112 27028 46121
rect 29644 46112 29696 46164
rect 33232 46155 33284 46164
rect 33232 46121 33241 46155
rect 33241 46121 33275 46155
rect 33275 46121 33284 46155
rect 33232 46112 33284 46121
rect 39948 46112 40000 46164
rect 45560 46112 45612 46164
rect 48044 46112 48096 46164
rect 14648 46044 14700 46096
rect 1768 46019 1820 46028
rect 1768 45985 1777 46019
rect 1777 45985 1811 46019
rect 1811 45985 1820 46019
rect 1768 45976 1820 45985
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 4896 46019 4948 46028
rect 4896 45985 4905 46019
rect 4905 45985 4939 46019
rect 4939 45985 4948 46019
rect 4896 45976 4948 45985
rect 5540 45976 5592 46028
rect 5816 45976 5868 46028
rect 10416 46019 10468 46028
rect 10416 45985 10425 46019
rect 10425 45985 10459 46019
rect 10459 45985 10468 46019
rect 10416 45976 10468 45985
rect 10968 45976 11020 46028
rect 14556 45976 14608 46028
rect 14832 46019 14884 46028
rect 14832 45985 14841 46019
rect 14841 45985 14875 46019
rect 14875 45985 14884 46019
rect 14832 45976 14884 45985
rect 4804 45908 4856 45960
rect 13360 45908 13412 45960
rect 13544 45951 13596 45960
rect 13544 45917 13553 45951
rect 13553 45917 13587 45951
rect 13587 45917 13596 45951
rect 13544 45908 13596 45917
rect 16580 45951 16632 45960
rect 16580 45917 16589 45951
rect 16589 45917 16623 45951
rect 16623 45917 16632 45951
rect 41512 46044 41564 46096
rect 45376 46044 45428 46096
rect 47032 46044 47084 46096
rect 25136 46019 25188 46028
rect 25136 45985 25145 46019
rect 25145 45985 25179 46019
rect 25179 45985 25188 46019
rect 25136 45976 25188 45985
rect 29920 45976 29972 46028
rect 30288 45976 30340 46028
rect 35532 46019 35584 46028
rect 35532 45985 35541 46019
rect 35541 45985 35575 46019
rect 35575 45985 35584 46019
rect 35532 45976 35584 45985
rect 36084 46019 36136 46028
rect 36084 45985 36093 46019
rect 36093 45985 36127 46019
rect 36127 45985 36136 46019
rect 36084 45976 36136 45985
rect 40592 46019 40644 46028
rect 40592 45985 40601 46019
rect 40601 45985 40635 46019
rect 40635 45985 40644 46019
rect 40592 45976 40644 45985
rect 45744 46019 45796 46028
rect 45744 45985 45753 46019
rect 45753 45985 45787 46019
rect 45787 45985 45796 46019
rect 45744 45976 45796 45985
rect 16580 45908 16632 45917
rect 3056 45840 3108 45892
rect 6644 45840 6696 45892
rect 10600 45883 10652 45892
rect 10600 45849 10609 45883
rect 10609 45849 10643 45883
rect 10643 45849 10652 45883
rect 10600 45840 10652 45849
rect 26976 45908 27028 45960
rect 29000 45951 29052 45960
rect 29000 45917 29009 45951
rect 29009 45917 29043 45951
rect 29043 45917 29052 45951
rect 29000 45908 29052 45917
rect 37924 45951 37976 45960
rect 24768 45883 24820 45892
rect 24768 45849 24777 45883
rect 24777 45849 24811 45883
rect 24811 45849 24820 45883
rect 24768 45840 24820 45849
rect 29920 45883 29972 45892
rect 29920 45849 29929 45883
rect 29929 45849 29963 45883
rect 29963 45849 29972 45883
rect 29920 45840 29972 45849
rect 22836 45772 22888 45824
rect 37924 45917 37933 45951
rect 37933 45917 37967 45951
rect 37967 45917 37976 45951
rect 37924 45908 37976 45917
rect 40132 45951 40184 45960
rect 40132 45917 40141 45951
rect 40141 45917 40175 45951
rect 40175 45917 40184 45951
rect 40132 45908 40184 45917
rect 35716 45883 35768 45892
rect 35716 45849 35725 45883
rect 35725 45849 35759 45883
rect 35759 45849 35768 45883
rect 35716 45840 35768 45849
rect 40316 45883 40368 45892
rect 40316 45849 40325 45883
rect 40325 45849 40359 45883
rect 40359 45849 40368 45883
rect 40316 45840 40368 45849
rect 45928 45883 45980 45892
rect 45928 45849 45937 45883
rect 45937 45849 45971 45883
rect 45971 45849 45980 45883
rect 45928 45840 45980 45849
rect 47584 45772 47636 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 6644 45611 6696 45620
rect 6644 45577 6653 45611
rect 6653 45577 6687 45611
rect 6687 45577 6696 45611
rect 6644 45568 6696 45577
rect 10600 45611 10652 45620
rect 10600 45577 10609 45611
rect 10609 45577 10643 45611
rect 10643 45577 10652 45611
rect 10600 45568 10652 45577
rect 13544 45568 13596 45620
rect 12440 45543 12492 45552
rect 12440 45509 12449 45543
rect 12449 45509 12483 45543
rect 12483 45509 12492 45543
rect 12440 45500 12492 45509
rect 4712 45475 4764 45484
rect 4712 45441 4721 45475
rect 4721 45441 4755 45475
rect 4755 45441 4764 45475
rect 4712 45432 4764 45441
rect 4896 45432 4948 45484
rect 2504 45364 2556 45416
rect 2964 45407 3016 45416
rect 2964 45373 2973 45407
rect 2973 45373 3007 45407
rect 3007 45373 3016 45407
rect 2964 45364 3016 45373
rect 4988 45407 5040 45416
rect 4988 45373 4997 45407
rect 4997 45373 5031 45407
rect 5031 45373 5040 45407
rect 4988 45364 5040 45373
rect 10324 45364 10376 45416
rect 2320 45296 2372 45348
rect 10508 45475 10560 45484
rect 10508 45441 10517 45475
rect 10517 45441 10551 45475
rect 10551 45441 10560 45475
rect 12348 45475 12400 45484
rect 10508 45432 10560 45441
rect 12348 45441 12357 45475
rect 12357 45441 12391 45475
rect 12391 45441 12400 45475
rect 12348 45432 12400 45441
rect 12992 45475 13044 45484
rect 12992 45441 13001 45475
rect 13001 45441 13035 45475
rect 13035 45441 13044 45475
rect 12992 45432 13044 45441
rect 13360 45432 13412 45484
rect 24768 45568 24820 45620
rect 24952 45568 25004 45620
rect 29920 45568 29972 45620
rect 35716 45611 35768 45620
rect 29000 45500 29052 45552
rect 29736 45475 29788 45484
rect 29736 45441 29745 45475
rect 29745 45441 29779 45475
rect 29779 45441 29788 45475
rect 29736 45432 29788 45441
rect 35716 45577 35725 45611
rect 35725 45577 35759 45611
rect 35759 45577 35768 45611
rect 35716 45568 35768 45577
rect 37648 45500 37700 45552
rect 42800 45500 42852 45552
rect 47860 45500 47912 45552
rect 35624 45475 35676 45484
rect 35624 45441 35633 45475
rect 35633 45441 35667 45475
rect 35667 45441 35676 45475
rect 35624 45432 35676 45441
rect 36544 45475 36596 45484
rect 36544 45441 36553 45475
rect 36553 45441 36587 45475
rect 36587 45441 36596 45475
rect 36544 45432 36596 45441
rect 37924 45432 37976 45484
rect 40132 45432 40184 45484
rect 41512 45475 41564 45484
rect 41512 45441 41521 45475
rect 41521 45441 41555 45475
rect 41555 45441 41564 45475
rect 41512 45432 41564 45441
rect 14188 45407 14240 45416
rect 14188 45373 14197 45407
rect 14197 45373 14231 45407
rect 14231 45373 14240 45407
rect 14188 45364 14240 45373
rect 46848 45407 46900 45416
rect 46848 45373 46857 45407
rect 46857 45373 46891 45407
rect 46891 45373 46900 45407
rect 46848 45364 46900 45373
rect 26976 45296 27028 45348
rect 2228 45228 2280 45280
rect 12348 45228 12400 45280
rect 16580 45228 16632 45280
rect 46480 45228 46532 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 4620 45024 4672 45076
rect 40316 45067 40368 45076
rect 40316 45033 40325 45067
rect 40325 45033 40359 45067
rect 40359 45033 40368 45067
rect 40316 45024 40368 45033
rect 45928 45024 45980 45076
rect 1768 44863 1820 44872
rect 1768 44829 1777 44863
rect 1777 44829 1811 44863
rect 1811 44829 1820 44863
rect 1768 44820 1820 44829
rect 2412 44684 2464 44736
rect 22836 44888 22888 44940
rect 46480 44931 46532 44940
rect 46480 44897 46489 44931
rect 46489 44897 46523 44931
rect 46523 44897 46532 44931
rect 46480 44888 46532 44897
rect 48228 44931 48280 44940
rect 48228 44897 48237 44931
rect 48237 44897 48271 44931
rect 48271 44897 48280 44931
rect 48228 44888 48280 44897
rect 4896 44820 4948 44872
rect 40224 44863 40276 44872
rect 3240 44795 3292 44804
rect 3240 44761 3249 44795
rect 3249 44761 3283 44795
rect 3283 44761 3292 44795
rect 3240 44752 3292 44761
rect 40224 44829 40233 44863
rect 40233 44829 40267 44863
rect 40267 44829 40276 44863
rect 40224 44820 40276 44829
rect 4528 44684 4580 44736
rect 4712 44684 4764 44736
rect 5724 44752 5776 44804
rect 12348 44752 12400 44804
rect 46664 44795 46716 44804
rect 46664 44761 46673 44795
rect 46673 44761 46707 44795
rect 46707 44761 46716 44795
rect 46664 44752 46716 44761
rect 47676 44684 47728 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 2504 44480 2556 44532
rect 46664 44480 46716 44532
rect 2412 44455 2464 44464
rect 2412 44421 2421 44455
rect 2421 44421 2455 44455
rect 2455 44421 2464 44455
rect 2412 44412 2464 44421
rect 7380 44455 7432 44464
rect 7380 44421 7389 44455
rect 7389 44421 7423 44455
rect 7423 44421 7432 44455
rect 7380 44412 7432 44421
rect 12992 44412 13044 44464
rect 2228 44387 2280 44396
rect 2228 44353 2237 44387
rect 2237 44353 2271 44387
rect 2271 44353 2280 44387
rect 2228 44344 2280 44353
rect 4528 44387 4580 44396
rect 4528 44353 4537 44387
rect 4537 44353 4571 44387
rect 4571 44353 4580 44387
rect 4528 44344 4580 44353
rect 2780 44319 2832 44328
rect 2780 44285 2789 44319
rect 2789 44285 2823 44319
rect 2823 44285 2832 44319
rect 2780 44276 2832 44285
rect 5448 44319 5500 44328
rect 5448 44285 5457 44319
rect 5457 44285 5491 44319
rect 5491 44285 5500 44319
rect 41512 44344 41564 44396
rect 47768 44344 47820 44396
rect 48320 44387 48372 44396
rect 48320 44353 48329 44387
rect 48329 44353 48363 44387
rect 48363 44353 48372 44387
rect 48320 44344 48372 44353
rect 5448 44276 5500 44285
rect 40224 44276 40276 44328
rect 3976 44208 4028 44260
rect 47216 44183 47268 44192
rect 47216 44149 47225 44183
rect 47225 44149 47259 44183
rect 47259 44149 47268 44183
rect 47216 44140 47268 44149
rect 47308 44140 47360 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 4068 43979 4120 43988
rect 4068 43945 4077 43979
rect 4077 43945 4111 43979
rect 4111 43945 4120 43979
rect 4068 43936 4120 43945
rect 2780 43843 2832 43852
rect 2780 43809 2789 43843
rect 2789 43809 2823 43843
rect 2823 43809 2832 43843
rect 2780 43800 2832 43809
rect 4988 43800 5040 43852
rect 5540 43843 5592 43852
rect 5540 43809 5549 43843
rect 5549 43809 5583 43843
rect 5583 43809 5592 43843
rect 5540 43800 5592 43809
rect 47216 43800 47268 43852
rect 48136 43843 48188 43852
rect 48136 43809 48145 43843
rect 48145 43809 48179 43843
rect 48179 43809 48188 43843
rect 48136 43800 48188 43809
rect 1584 43775 1636 43784
rect 1584 43741 1593 43775
rect 1593 43741 1627 43775
rect 1627 43741 1636 43775
rect 1584 43732 1636 43741
rect 3976 43775 4028 43784
rect 3976 43741 3985 43775
rect 3985 43741 4019 43775
rect 4019 43741 4028 43775
rect 3976 43732 4028 43741
rect 4712 43732 4764 43784
rect 2596 43664 2648 43716
rect 5540 43664 5592 43716
rect 13544 43664 13596 43716
rect 27804 43732 27856 43784
rect 27436 43664 27488 43716
rect 47124 43664 47176 43716
rect 27344 43639 27396 43648
rect 27344 43605 27353 43639
rect 27353 43605 27387 43639
rect 27387 43605 27396 43639
rect 27344 43596 27396 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 2596 43435 2648 43444
rect 2596 43401 2605 43435
rect 2605 43401 2639 43435
rect 2639 43401 2648 43435
rect 2596 43392 2648 43401
rect 4620 43392 4672 43444
rect 47124 43435 47176 43444
rect 7840 43324 7892 43376
rect 22376 43324 22428 43376
rect 1584 43256 1636 43308
rect 1952 43188 2004 43240
rect 4712 43256 4764 43308
rect 9128 43256 9180 43308
rect 4620 43231 4672 43240
rect 4620 43197 4629 43231
rect 4629 43197 4663 43231
rect 4663 43197 4672 43231
rect 4620 43188 4672 43197
rect 22560 43256 22612 43308
rect 29736 43324 29788 43376
rect 27344 43299 27396 43308
rect 27344 43265 27353 43299
rect 27353 43265 27387 43299
rect 27387 43265 27396 43299
rect 27344 43256 27396 43265
rect 28540 43256 28592 43308
rect 29000 43256 29052 43308
rect 30472 43299 30524 43308
rect 30472 43265 30481 43299
rect 30481 43265 30515 43299
rect 30515 43265 30524 43299
rect 30472 43256 30524 43265
rect 36084 43256 36136 43308
rect 27436 43188 27488 43240
rect 47124 43401 47133 43435
rect 47133 43401 47167 43435
rect 47167 43401 47176 43435
rect 47124 43392 47176 43401
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 47492 43256 47544 43308
rect 23664 43120 23716 43172
rect 23572 43052 23624 43104
rect 27252 43052 27304 43104
rect 29828 43095 29880 43104
rect 29828 43061 29837 43095
rect 29837 43061 29871 43095
rect 29871 43061 29880 43095
rect 29828 43052 29880 43061
rect 30288 43095 30340 43104
rect 30288 43061 30297 43095
rect 30297 43061 30331 43095
rect 30331 43061 30340 43095
rect 30288 43052 30340 43061
rect 35900 43052 35952 43104
rect 47860 43095 47912 43104
rect 47860 43061 47869 43095
rect 47869 43061 47903 43095
rect 47903 43061 47912 43095
rect 47860 43052 47912 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 2320 42712 2372 42764
rect 3056 42755 3108 42764
rect 3056 42721 3065 42755
rect 3065 42721 3099 42755
rect 3099 42721 3108 42755
rect 3056 42712 3108 42721
rect 4712 42755 4764 42764
rect 4712 42721 4721 42755
rect 4721 42721 4755 42755
rect 4755 42721 4764 42755
rect 4712 42712 4764 42721
rect 28080 42712 28132 42764
rect 28540 42712 28592 42764
rect 47860 42712 47912 42764
rect 48228 42755 48280 42764
rect 48228 42721 48237 42755
rect 48237 42721 48271 42755
rect 48271 42721 48280 42755
rect 48228 42712 48280 42721
rect 2872 42644 2924 42696
rect 4804 42644 4856 42696
rect 23664 42687 23716 42696
rect 23664 42653 23673 42687
rect 23673 42653 23707 42687
rect 23707 42653 23716 42687
rect 23664 42644 23716 42653
rect 28448 42687 28500 42696
rect 28448 42653 28457 42687
rect 28457 42653 28491 42687
rect 28491 42653 28500 42687
rect 28448 42644 28500 42653
rect 28724 42644 28776 42696
rect 30288 42644 30340 42696
rect 32128 42644 32180 42696
rect 35348 42644 35400 42696
rect 28908 42576 28960 42628
rect 32864 42576 32916 42628
rect 33876 42576 33928 42628
rect 35900 42644 35952 42696
rect 2688 42508 2740 42560
rect 23480 42551 23532 42560
rect 23480 42517 23489 42551
rect 23489 42517 23523 42551
rect 23523 42517 23532 42551
rect 23480 42508 23532 42517
rect 27344 42551 27396 42560
rect 27344 42517 27353 42551
rect 27353 42517 27387 42551
rect 27387 42517 27396 42551
rect 27344 42508 27396 42517
rect 29184 42508 29236 42560
rect 31116 42551 31168 42560
rect 31116 42517 31125 42551
rect 31125 42517 31159 42551
rect 31159 42517 31168 42551
rect 31116 42508 31168 42517
rect 32404 42508 32456 42560
rect 34888 42551 34940 42560
rect 34888 42517 34897 42551
rect 34897 42517 34931 42551
rect 34931 42517 34940 42551
rect 34888 42508 34940 42517
rect 37188 42551 37240 42560
rect 37188 42517 37197 42551
rect 37197 42517 37231 42551
rect 37231 42517 37240 42551
rect 37188 42508 37240 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 4712 42236 4764 42288
rect 23480 42236 23532 42288
rect 23572 42211 23624 42220
rect 23572 42177 23581 42211
rect 23581 42177 23615 42211
rect 23615 42177 23624 42211
rect 23572 42168 23624 42177
rect 24308 42168 24360 42220
rect 28080 42236 28132 42288
rect 28724 42236 28776 42288
rect 27252 42168 27304 42220
rect 29184 42211 29236 42220
rect 29184 42177 29193 42211
rect 29193 42177 29227 42211
rect 29227 42177 29236 42211
rect 29184 42168 29236 42177
rect 29828 42211 29880 42220
rect 29828 42177 29837 42211
rect 29837 42177 29871 42211
rect 29871 42177 29880 42211
rect 29828 42168 29880 42177
rect 30472 42236 30524 42288
rect 32864 42304 32916 42356
rect 36084 42347 36136 42356
rect 36084 42313 36093 42347
rect 36093 42313 36127 42347
rect 36127 42313 36136 42347
rect 36084 42304 36136 42313
rect 31116 42211 31168 42220
rect 31116 42177 31125 42211
rect 31125 42177 31159 42211
rect 31159 42177 31168 42211
rect 31116 42168 31168 42177
rect 36544 42236 36596 42288
rect 32496 42211 32548 42220
rect 30564 42100 30616 42152
rect 29000 42075 29052 42084
rect 29000 42041 29009 42075
rect 29009 42041 29043 42075
rect 29043 42041 29052 42075
rect 29000 42032 29052 42041
rect 32496 42177 32505 42211
rect 32505 42177 32539 42211
rect 32539 42177 32548 42211
rect 32496 42168 32548 42177
rect 33876 42211 33928 42220
rect 33876 42177 33885 42211
rect 33885 42177 33919 42211
rect 33919 42177 33928 42211
rect 33876 42168 33928 42177
rect 34888 42168 34940 42220
rect 35900 42211 35952 42220
rect 35900 42177 35909 42211
rect 35909 42177 35943 42211
rect 35943 42177 35952 42211
rect 35900 42168 35952 42177
rect 37648 42211 37700 42220
rect 37648 42177 37657 42211
rect 37657 42177 37691 42211
rect 37691 42177 37700 42211
rect 37648 42168 37700 42177
rect 38568 42168 38620 42220
rect 47308 42236 47360 42288
rect 43444 42168 43496 42220
rect 47768 42211 47820 42220
rect 47768 42177 47777 42211
rect 47777 42177 47811 42211
rect 47811 42177 47820 42211
rect 47768 42168 47820 42177
rect 33140 42032 33192 42084
rect 37188 42100 37240 42152
rect 38752 42100 38804 42152
rect 42616 42143 42668 42152
rect 42616 42109 42625 42143
rect 42625 42109 42659 42143
rect 42659 42109 42668 42143
rect 42616 42100 42668 42109
rect 23388 42007 23440 42016
rect 23388 41973 23397 42007
rect 23397 41973 23431 42007
rect 23431 41973 23440 42007
rect 23388 41964 23440 41973
rect 27896 41964 27948 42016
rect 28540 42007 28592 42016
rect 28540 41973 28549 42007
rect 28549 41973 28583 42007
rect 28583 41973 28592 42007
rect 28540 41964 28592 41973
rect 32312 42007 32364 42016
rect 32312 41973 32321 42007
rect 32321 41973 32355 42007
rect 32355 41973 32364 42007
rect 32312 41964 32364 41973
rect 35532 41964 35584 42016
rect 36728 42007 36780 42016
rect 36728 41973 36737 42007
rect 36737 41973 36771 42007
rect 36771 41973 36780 42007
rect 36728 41964 36780 41973
rect 38292 42007 38344 42016
rect 38292 41973 38301 42007
rect 38301 41973 38335 42007
rect 38335 41973 38344 42007
rect 38292 41964 38344 41973
rect 40224 42007 40276 42016
rect 40224 41973 40233 42007
rect 40233 41973 40267 42007
rect 40267 41973 40276 42007
rect 40224 41964 40276 41973
rect 43996 42007 44048 42016
rect 43996 41973 44005 42007
rect 44005 41973 44039 42007
rect 44039 41973 44048 42007
rect 43996 41964 44048 41973
rect 46480 41964 46532 42016
rect 47860 42007 47912 42016
rect 47860 41973 47869 42007
rect 47869 41973 47903 42007
rect 47903 41973 47912 42007
rect 47860 41964 47912 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 28448 41760 28500 41812
rect 28632 41760 28684 41812
rect 28908 41803 28960 41812
rect 28908 41769 28917 41803
rect 28917 41769 28951 41803
rect 28951 41769 28960 41803
rect 28908 41760 28960 41769
rect 35348 41760 35400 41812
rect 35900 41760 35952 41812
rect 37648 41760 37700 41812
rect 38568 41803 38620 41812
rect 38568 41769 38577 41803
rect 38577 41769 38611 41803
rect 38611 41769 38620 41803
rect 38568 41760 38620 41769
rect 43444 41760 43496 41812
rect 31116 41692 31168 41744
rect 31484 41624 31536 41676
rect 2044 41556 2096 41608
rect 24308 41556 24360 41608
rect 28080 41556 28132 41608
rect 23388 41488 23440 41540
rect 27344 41488 27396 41540
rect 28724 41599 28776 41608
rect 28724 41565 28733 41599
rect 28733 41565 28767 41599
rect 28767 41565 28776 41599
rect 28724 41556 28776 41565
rect 30564 41556 30616 41608
rect 29920 41488 29972 41540
rect 30656 41488 30708 41540
rect 31024 41488 31076 41540
rect 30932 41463 30984 41472
rect 30932 41429 30941 41463
rect 30941 41429 30975 41463
rect 30975 41429 30984 41463
rect 32128 41556 32180 41608
rect 34796 41556 34848 41608
rect 38200 41667 38252 41676
rect 38200 41633 38209 41667
rect 38209 41633 38243 41667
rect 38243 41633 38252 41667
rect 38200 41624 38252 41633
rect 32312 41488 32364 41540
rect 34060 41488 34112 41540
rect 37464 41556 37516 41608
rect 37648 41556 37700 41608
rect 43168 41624 43220 41676
rect 46480 41667 46532 41676
rect 46480 41633 46489 41667
rect 46489 41633 46523 41667
rect 46523 41633 46532 41667
rect 46480 41624 46532 41633
rect 47860 41624 47912 41676
rect 48228 41667 48280 41676
rect 48228 41633 48237 41667
rect 48237 41633 48271 41667
rect 48271 41633 48280 41667
rect 48228 41624 48280 41633
rect 42892 41599 42944 41608
rect 42892 41565 42901 41599
rect 42901 41565 42935 41599
rect 42935 41565 42944 41599
rect 42892 41556 42944 41565
rect 36728 41488 36780 41540
rect 45560 41556 45612 41608
rect 44088 41488 44140 41540
rect 30932 41420 30984 41429
rect 37740 41463 37792 41472
rect 37740 41429 37749 41463
rect 37749 41429 37783 41463
rect 37783 41429 37792 41463
rect 37740 41420 37792 41429
rect 38200 41420 38252 41472
rect 45192 41463 45244 41472
rect 45192 41429 45201 41463
rect 45201 41429 45235 41463
rect 45235 41429 45244 41463
rect 45192 41420 45244 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 32496 41216 32548 41268
rect 33140 41216 33192 41268
rect 34060 41216 34112 41268
rect 35624 41216 35676 41268
rect 30932 41148 30984 41200
rect 2044 41123 2096 41132
rect 2044 41089 2053 41123
rect 2053 41089 2087 41123
rect 2087 41089 2096 41123
rect 2044 41080 2096 41089
rect 24308 41080 24360 41132
rect 24492 41123 24544 41132
rect 24492 41089 24526 41123
rect 24526 41089 24544 41123
rect 24492 41080 24544 41089
rect 31116 41080 31168 41132
rect 32404 41123 32456 41132
rect 32404 41089 32413 41123
rect 32413 41089 32447 41123
rect 32447 41089 32456 41123
rect 32404 41080 32456 41089
rect 37372 41148 37424 41200
rect 33968 41123 34020 41132
rect 33968 41089 33977 41123
rect 33977 41089 34011 41123
rect 34011 41089 34020 41123
rect 33968 41080 34020 41089
rect 2412 41012 2464 41064
rect 2780 41055 2832 41064
rect 2780 41021 2789 41055
rect 2789 41021 2823 41055
rect 2823 41021 2832 41055
rect 2780 41012 2832 41021
rect 30656 41055 30708 41064
rect 30656 41021 30665 41055
rect 30665 41021 30699 41055
rect 30699 41021 30708 41055
rect 30656 41012 30708 41021
rect 36544 41055 36596 41064
rect 36544 41021 36553 41055
rect 36553 41021 36587 41055
rect 36587 41021 36596 41055
rect 36544 41012 36596 41021
rect 37280 41080 37332 41132
rect 37740 41080 37792 41132
rect 38292 41148 38344 41200
rect 40224 41123 40276 41132
rect 37372 41012 37424 41064
rect 37464 41012 37516 41064
rect 25596 40919 25648 40928
rect 25596 40885 25605 40919
rect 25605 40885 25639 40919
rect 25639 40885 25648 40919
rect 25596 40876 25648 40885
rect 30564 40919 30616 40928
rect 30564 40885 30573 40919
rect 30573 40885 30607 40919
rect 30607 40885 30616 40919
rect 30564 40876 30616 40885
rect 30840 40876 30892 40928
rect 33784 40919 33836 40928
rect 33784 40885 33793 40919
rect 33793 40885 33827 40919
rect 33827 40885 33836 40919
rect 33784 40876 33836 40885
rect 37188 40944 37240 40996
rect 36636 40876 36688 40928
rect 40224 41089 40233 41123
rect 40233 41089 40267 41123
rect 40267 41089 40276 41123
rect 40224 41080 40276 41089
rect 41788 41080 41840 41132
rect 42892 41148 42944 41200
rect 45192 41148 45244 41200
rect 42248 41012 42300 41064
rect 43076 41123 43128 41132
rect 43076 41089 43085 41123
rect 43085 41089 43119 41123
rect 43119 41089 43128 41123
rect 43076 41080 43128 41089
rect 43996 41080 44048 41132
rect 44732 41080 44784 41132
rect 42892 41055 42944 41064
rect 42892 41021 42901 41055
rect 42901 41021 42935 41055
rect 42935 41021 42944 41055
rect 42892 41012 42944 41021
rect 39580 40987 39632 40996
rect 39580 40953 39589 40987
rect 39589 40953 39623 40987
rect 39623 40953 39632 40987
rect 39580 40944 39632 40953
rect 38568 40876 38620 40928
rect 39672 40876 39724 40928
rect 41144 40876 41196 40928
rect 42524 40876 42576 40928
rect 43168 40944 43220 40996
rect 43260 40919 43312 40928
rect 43260 40885 43269 40919
rect 43269 40885 43303 40919
rect 43303 40885 43312 40919
rect 43260 40876 43312 40885
rect 46480 40876 46532 40928
rect 47860 40919 47912 40928
rect 47860 40885 47869 40919
rect 47869 40885 47903 40919
rect 47903 40885 47912 40919
rect 47860 40876 47912 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 2412 40715 2464 40724
rect 2412 40681 2421 40715
rect 2421 40681 2455 40715
rect 2455 40681 2464 40715
rect 2412 40672 2464 40681
rect 24492 40672 24544 40724
rect 28264 40672 28316 40724
rect 28540 40715 28592 40724
rect 28540 40681 28549 40715
rect 28549 40681 28583 40715
rect 28583 40681 28592 40715
rect 28540 40672 28592 40681
rect 29920 40715 29972 40724
rect 29920 40681 29929 40715
rect 29929 40681 29963 40715
rect 29963 40681 29972 40715
rect 29920 40672 29972 40681
rect 34796 40672 34848 40724
rect 35808 40672 35860 40724
rect 42248 40715 42300 40724
rect 42248 40681 42257 40715
rect 42257 40681 42291 40715
rect 42291 40681 42300 40715
rect 42248 40672 42300 40681
rect 45560 40715 45612 40724
rect 45560 40681 45569 40715
rect 45569 40681 45603 40715
rect 45603 40681 45612 40715
rect 45560 40672 45612 40681
rect 28632 40604 28684 40656
rect 37280 40604 37332 40656
rect 2228 40468 2280 40520
rect 4712 40468 4764 40520
rect 24768 40511 24820 40520
rect 24768 40477 24777 40511
rect 24777 40477 24811 40511
rect 24811 40477 24820 40511
rect 32128 40536 32180 40588
rect 32956 40579 33008 40588
rect 32956 40545 32965 40579
rect 32965 40545 32999 40579
rect 32999 40545 33008 40579
rect 32956 40536 33008 40545
rect 38568 40536 38620 40588
rect 44088 40536 44140 40588
rect 46480 40579 46532 40588
rect 24768 40468 24820 40477
rect 33784 40468 33836 40520
rect 25044 40400 25096 40452
rect 29736 40443 29788 40452
rect 29736 40409 29745 40443
rect 29745 40409 29779 40443
rect 29779 40409 29788 40443
rect 29736 40400 29788 40409
rect 31024 40400 31076 40452
rect 34520 40400 34572 40452
rect 37096 40443 37148 40452
rect 37096 40409 37105 40443
rect 37105 40409 37139 40443
rect 37139 40409 37148 40443
rect 37096 40400 37148 40409
rect 37372 40400 37424 40452
rect 39580 40468 39632 40520
rect 40224 40511 40276 40520
rect 40224 40477 40233 40511
rect 40233 40477 40267 40511
rect 40267 40477 40276 40511
rect 41144 40511 41196 40520
rect 40224 40468 40276 40477
rect 41144 40477 41178 40511
rect 41178 40477 41196 40511
rect 41144 40468 41196 40477
rect 42616 40468 42668 40520
rect 44732 40468 44784 40520
rect 45284 40511 45336 40520
rect 45284 40477 45293 40511
rect 45293 40477 45327 40511
rect 45327 40477 45336 40511
rect 45284 40468 45336 40477
rect 46480 40545 46489 40579
rect 46489 40545 46523 40579
rect 46523 40545 46532 40579
rect 46480 40536 46532 40545
rect 47860 40536 47912 40588
rect 48228 40579 48280 40588
rect 48228 40545 48237 40579
rect 48237 40545 48271 40579
rect 48271 40545 48280 40579
rect 48228 40536 48280 40545
rect 41604 40400 41656 40452
rect 42800 40400 42852 40452
rect 42984 40443 43036 40452
rect 42984 40409 43018 40443
rect 43018 40409 43036 40443
rect 42984 40400 43036 40409
rect 29828 40332 29880 40384
rect 30104 40375 30156 40384
rect 30104 40341 30113 40375
rect 30113 40341 30147 40375
rect 30147 40341 30156 40375
rect 30104 40332 30156 40341
rect 35348 40332 35400 40384
rect 36544 40332 36596 40384
rect 37188 40375 37240 40384
rect 37188 40341 37197 40375
rect 37197 40341 37231 40375
rect 37231 40341 37240 40375
rect 37188 40332 37240 40341
rect 39212 40375 39264 40384
rect 39212 40341 39221 40375
rect 39221 40341 39255 40375
rect 39255 40341 39264 40375
rect 39212 40332 39264 40341
rect 42892 40332 42944 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 25044 40171 25096 40180
rect 25044 40137 25053 40171
rect 25053 40137 25087 40171
rect 25087 40137 25096 40171
rect 25044 40128 25096 40137
rect 29920 40128 29972 40180
rect 34520 40171 34572 40180
rect 34520 40137 34529 40171
rect 34529 40137 34563 40171
rect 34563 40137 34572 40171
rect 34520 40128 34572 40137
rect 35808 40128 35860 40180
rect 23940 40035 23992 40044
rect 23940 40001 23974 40035
rect 23974 40001 23992 40035
rect 25596 40035 25648 40044
rect 23940 39992 23992 40001
rect 25596 40001 25605 40035
rect 25605 40001 25639 40035
rect 25639 40001 25648 40035
rect 25596 39992 25648 40001
rect 24768 39924 24820 39976
rect 24308 39788 24360 39840
rect 24584 39788 24636 39840
rect 26608 39788 26660 39840
rect 30012 39992 30064 40044
rect 30840 40035 30892 40044
rect 30840 40001 30849 40035
rect 30849 40001 30883 40035
rect 30883 40001 30892 40035
rect 30840 39992 30892 40001
rect 30932 40035 30984 40044
rect 30932 40001 30941 40035
rect 30941 40001 30975 40035
rect 30975 40001 30984 40035
rect 30932 39992 30984 40001
rect 32956 39992 33008 40044
rect 33232 39992 33284 40044
rect 28080 39924 28132 39976
rect 29828 39924 29880 39976
rect 35348 40060 35400 40112
rect 35532 40103 35584 40112
rect 35532 40069 35541 40103
rect 35541 40069 35575 40103
rect 35575 40069 35584 40103
rect 35532 40060 35584 40069
rect 37188 40128 37240 40180
rect 42892 40171 42944 40180
rect 42892 40137 42901 40171
rect 42901 40137 42935 40171
rect 42935 40137 42944 40171
rect 42892 40128 42944 40137
rect 45284 40128 45336 40180
rect 39212 40060 39264 40112
rect 42248 40060 42300 40112
rect 36636 40035 36688 40044
rect 36636 40001 36645 40035
rect 36645 40001 36679 40035
rect 36679 40001 36688 40035
rect 36636 39992 36688 40001
rect 36728 40035 36780 40044
rect 36728 40001 36737 40035
rect 36737 40001 36771 40035
rect 36771 40001 36780 40035
rect 41604 40035 41656 40044
rect 36728 39992 36780 40001
rect 41604 40001 41613 40035
rect 41613 40001 41647 40035
rect 41647 40001 41656 40035
rect 41604 39992 41656 40001
rect 41788 40035 41840 40044
rect 41788 40001 41797 40035
rect 41797 40001 41831 40035
rect 41831 40001 41840 40035
rect 41788 39992 41840 40001
rect 43168 40060 43220 40112
rect 44088 40035 44140 40044
rect 44088 40001 44097 40035
rect 44097 40001 44131 40035
rect 44131 40001 44140 40035
rect 44088 39992 44140 40001
rect 45008 40035 45060 40044
rect 45008 40001 45042 40035
rect 45042 40001 45060 40035
rect 47768 40035 47820 40044
rect 45008 39992 45060 40001
rect 47768 40001 47777 40035
rect 47777 40001 47811 40035
rect 47811 40001 47820 40035
rect 47768 39992 47820 40001
rect 35808 39967 35860 39976
rect 35808 39933 35817 39967
rect 35817 39933 35851 39967
rect 35851 39933 35860 39967
rect 35808 39924 35860 39933
rect 38108 39924 38160 39976
rect 38568 39924 38620 39976
rect 43076 39924 43128 39976
rect 44180 39924 44232 39976
rect 44732 39967 44784 39976
rect 44732 39933 44741 39967
rect 44741 39933 44775 39967
rect 44775 39933 44784 39967
rect 44732 39924 44784 39933
rect 30380 39856 30432 39908
rect 35440 39856 35492 39908
rect 30472 39831 30524 39840
rect 30472 39797 30481 39831
rect 30481 39797 30515 39831
rect 30515 39797 30524 39831
rect 30472 39788 30524 39797
rect 35716 39788 35768 39840
rect 42800 39788 42852 39840
rect 45376 39788 45428 39840
rect 46480 39788 46532 39840
rect 47860 39831 47912 39840
rect 47860 39797 47869 39831
rect 47869 39797 47903 39831
rect 47903 39797 47912 39831
rect 47860 39788 47912 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 23940 39584 23992 39636
rect 30012 39584 30064 39636
rect 33232 39584 33284 39636
rect 33968 39584 34020 39636
rect 35440 39627 35492 39636
rect 24584 39516 24636 39568
rect 35440 39593 35449 39627
rect 35449 39593 35483 39627
rect 35483 39593 35492 39627
rect 35440 39584 35492 39593
rect 42984 39584 43036 39636
rect 45008 39584 45060 39636
rect 24768 39423 24820 39432
rect 24768 39389 24777 39423
rect 24777 39389 24811 39423
rect 24811 39389 24820 39423
rect 28264 39448 28316 39500
rect 24768 39380 24820 39389
rect 28172 39380 28224 39432
rect 30104 39448 30156 39500
rect 28632 39423 28684 39432
rect 28632 39389 28641 39423
rect 28641 39389 28675 39423
rect 28675 39389 28684 39423
rect 28632 39380 28684 39389
rect 28908 39423 28960 39432
rect 28908 39389 28917 39423
rect 28917 39389 28951 39423
rect 28951 39389 28960 39423
rect 28908 39380 28960 39389
rect 29736 39423 29788 39432
rect 29736 39389 29745 39423
rect 29745 39389 29779 39423
rect 29779 39389 29788 39423
rect 29736 39380 29788 39389
rect 30380 39380 30432 39432
rect 31300 39380 31352 39432
rect 31484 39380 31536 39432
rect 26424 39312 26476 39364
rect 28540 39355 28592 39364
rect 28540 39321 28549 39355
rect 28549 39321 28583 39355
rect 28583 39321 28592 39355
rect 28540 39312 28592 39321
rect 30472 39312 30524 39364
rect 32036 39380 32088 39432
rect 34060 39423 34112 39432
rect 34060 39389 34069 39423
rect 34069 39389 34103 39423
rect 34103 39389 34112 39423
rect 35532 39448 35584 39500
rect 46480 39491 46532 39500
rect 46480 39457 46489 39491
rect 46489 39457 46523 39491
rect 46523 39457 46532 39491
rect 46480 39448 46532 39457
rect 47860 39448 47912 39500
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 34060 39380 34112 39389
rect 38108 39423 38160 39432
rect 34520 39312 34572 39364
rect 38108 39389 38117 39423
rect 38117 39389 38151 39423
rect 38151 39389 38160 39423
rect 38108 39380 38160 39389
rect 39672 39380 39724 39432
rect 42524 39423 42576 39432
rect 42524 39389 42533 39423
rect 42533 39389 42567 39423
rect 42567 39389 42576 39423
rect 42524 39380 42576 39389
rect 45376 39423 45428 39432
rect 45376 39389 45385 39423
rect 45385 39389 45419 39423
rect 45419 39389 45428 39423
rect 45376 39380 45428 39389
rect 37556 39312 37608 39364
rect 25596 39244 25648 39296
rect 25688 39244 25740 39296
rect 27804 39287 27856 39296
rect 27804 39253 27813 39287
rect 27813 39253 27847 39287
rect 27847 39253 27856 39287
rect 27804 39244 27856 39253
rect 28356 39244 28408 39296
rect 34060 39244 34112 39296
rect 38660 39244 38712 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 25688 39083 25740 39092
rect 25688 39049 25697 39083
rect 25697 39049 25731 39083
rect 25731 39049 25740 39083
rect 25688 39040 25740 39049
rect 25780 39083 25832 39092
rect 25780 39049 25789 39083
rect 25789 39049 25823 39083
rect 25823 39049 25832 39083
rect 26424 39083 26476 39092
rect 25780 39040 25832 39049
rect 26424 39049 26433 39083
rect 26433 39049 26467 39083
rect 26467 39049 26476 39083
rect 26424 39040 26476 39049
rect 29736 39040 29788 39092
rect 25044 38972 25096 39024
rect 25596 39015 25648 39024
rect 25596 38981 25605 39015
rect 25605 38981 25639 39015
rect 25639 38981 25648 39015
rect 25596 38972 25648 38981
rect 28540 38972 28592 39024
rect 28908 38972 28960 39024
rect 26608 38947 26660 38956
rect 26608 38913 26617 38947
rect 26617 38913 26651 38947
rect 26651 38913 26660 38947
rect 26608 38904 26660 38913
rect 28080 38947 28132 38956
rect 28080 38913 28089 38947
rect 28089 38913 28123 38947
rect 28123 38913 28132 38947
rect 28080 38904 28132 38913
rect 31208 38947 31260 38956
rect 31208 38913 31217 38947
rect 31217 38913 31251 38947
rect 31251 38913 31260 38947
rect 31208 38904 31260 38913
rect 32036 38904 32088 38956
rect 36728 39040 36780 39092
rect 40224 39040 40276 39092
rect 35716 39015 35768 39024
rect 35716 38981 35750 39015
rect 35750 38981 35768 39015
rect 35716 38972 35768 38981
rect 43260 38972 43312 39024
rect 37556 38904 37608 38956
rect 39028 38904 39080 38956
rect 44180 38947 44232 38956
rect 44180 38913 44189 38947
rect 44189 38913 44223 38947
rect 44223 38913 44232 38947
rect 44180 38904 44232 38913
rect 44456 38947 44508 38956
rect 44456 38913 44465 38947
rect 44465 38913 44499 38947
rect 44499 38913 44508 38947
rect 44456 38904 44508 38913
rect 45560 38904 45612 38956
rect 33048 38836 33100 38888
rect 25964 38743 26016 38752
rect 25964 38709 25973 38743
rect 25973 38709 26007 38743
rect 26007 38709 26016 38743
rect 25964 38700 26016 38709
rect 31116 38700 31168 38752
rect 31300 38700 31352 38752
rect 34612 38768 34664 38820
rect 32864 38700 32916 38752
rect 35808 38700 35860 38752
rect 43536 38836 43588 38888
rect 44364 38879 44416 38888
rect 44364 38845 44373 38879
rect 44373 38845 44407 38879
rect 44407 38845 44416 38879
rect 44364 38836 44416 38845
rect 45284 38836 45336 38888
rect 45468 38836 45520 38888
rect 43720 38743 43772 38752
rect 43720 38709 43729 38743
rect 43729 38709 43763 38743
rect 43763 38709 43772 38743
rect 43720 38700 43772 38709
rect 44272 38743 44324 38752
rect 44272 38709 44281 38743
rect 44281 38709 44315 38743
rect 44315 38709 44324 38743
rect 44272 38700 44324 38709
rect 44548 38700 44600 38752
rect 47952 38743 48004 38752
rect 47952 38709 47961 38743
rect 47961 38709 47995 38743
rect 47995 38709 48004 38743
rect 47952 38700 48004 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 25596 38539 25648 38548
rect 25596 38505 25605 38539
rect 25605 38505 25639 38539
rect 25639 38505 25648 38539
rect 25596 38496 25648 38505
rect 28540 38539 28592 38548
rect 28540 38505 28549 38539
rect 28549 38505 28583 38539
rect 28583 38505 28592 38539
rect 28540 38496 28592 38505
rect 25688 38403 25740 38412
rect 25688 38369 25697 38403
rect 25697 38369 25731 38403
rect 25731 38369 25740 38403
rect 25688 38360 25740 38369
rect 32128 38496 32180 38548
rect 40040 38539 40092 38548
rect 40040 38505 40049 38539
rect 40049 38505 40083 38539
rect 40083 38505 40092 38539
rect 45560 38539 45612 38548
rect 40040 38496 40092 38505
rect 33416 38360 33468 38412
rect 36728 38360 36780 38412
rect 37188 38360 37240 38412
rect 24768 38335 24820 38344
rect 24768 38301 24777 38335
rect 24777 38301 24811 38335
rect 24811 38301 24820 38335
rect 24768 38292 24820 38301
rect 25044 38292 25096 38344
rect 27804 38292 27856 38344
rect 31116 38335 31168 38344
rect 31116 38301 31150 38335
rect 31150 38301 31168 38335
rect 31116 38292 31168 38301
rect 32864 38335 32916 38344
rect 32864 38301 32873 38335
rect 32873 38301 32907 38335
rect 32907 38301 32916 38335
rect 32864 38292 32916 38301
rect 37096 38335 37148 38344
rect 37096 38301 37105 38335
rect 37105 38301 37139 38335
rect 37139 38301 37148 38335
rect 37096 38292 37148 38301
rect 38752 38292 38804 38344
rect 25688 38224 25740 38276
rect 39028 38335 39080 38344
rect 39028 38301 39037 38335
rect 39037 38301 39071 38335
rect 39071 38301 39080 38335
rect 39028 38292 39080 38301
rect 43076 38360 43128 38412
rect 23848 38156 23900 38208
rect 26240 38156 26292 38208
rect 33508 38199 33560 38208
rect 33508 38165 33517 38199
rect 33517 38165 33551 38199
rect 33551 38165 33560 38199
rect 33508 38156 33560 38165
rect 36912 38156 36964 38208
rect 39948 38156 40000 38208
rect 42800 38335 42852 38344
rect 42800 38301 42809 38335
rect 42809 38301 42843 38335
rect 42843 38301 42852 38335
rect 45560 38505 45569 38539
rect 45569 38505 45603 38539
rect 45603 38505 45612 38539
rect 45560 38496 45612 38505
rect 44456 38428 44508 38480
rect 45100 38428 45152 38480
rect 43352 38360 43404 38412
rect 44732 38360 44784 38412
rect 45468 38360 45520 38412
rect 48044 38403 48096 38412
rect 48044 38369 48053 38403
rect 48053 38369 48087 38403
rect 48087 38369 48096 38403
rect 48044 38360 48096 38369
rect 42800 38292 42852 38301
rect 44272 38335 44324 38344
rect 44272 38301 44281 38335
rect 44281 38301 44315 38335
rect 44315 38301 44324 38335
rect 44272 38292 44324 38301
rect 44364 38335 44416 38344
rect 44364 38301 44373 38335
rect 44373 38301 44407 38335
rect 44407 38301 44416 38335
rect 44364 38292 44416 38301
rect 45100 38292 45152 38344
rect 45376 38335 45428 38344
rect 45376 38301 45385 38335
rect 45385 38301 45419 38335
rect 45419 38301 45428 38335
rect 45376 38292 45428 38301
rect 46112 38292 46164 38344
rect 42892 38267 42944 38276
rect 42892 38233 42901 38267
rect 42901 38233 42935 38267
rect 42935 38233 42944 38267
rect 42892 38224 42944 38233
rect 43720 38224 43772 38276
rect 46848 38224 46900 38276
rect 44548 38156 44600 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 25596 37952 25648 38004
rect 29460 37995 29512 38004
rect 29460 37961 29469 37995
rect 29469 37961 29503 37995
rect 29503 37961 29512 37995
rect 29460 37952 29512 37961
rect 30932 37952 30984 38004
rect 31208 37952 31260 38004
rect 23848 37927 23900 37936
rect 23848 37893 23882 37927
rect 23882 37893 23900 37927
rect 23848 37884 23900 37893
rect 33508 37884 33560 37936
rect 24584 37816 24636 37868
rect 28080 37859 28132 37868
rect 28080 37825 28089 37859
rect 28089 37825 28123 37859
rect 28123 37825 28132 37859
rect 28080 37816 28132 37825
rect 28356 37859 28408 37868
rect 28356 37825 28390 37859
rect 28390 37825 28408 37859
rect 28356 37816 28408 37825
rect 31208 37859 31260 37868
rect 31208 37825 31217 37859
rect 31217 37825 31251 37859
rect 31251 37825 31260 37859
rect 31208 37816 31260 37825
rect 32128 37816 32180 37868
rect 36912 37859 36964 37868
rect 36912 37825 36921 37859
rect 36921 37825 36955 37859
rect 36955 37825 36964 37859
rect 36912 37816 36964 37825
rect 45100 37995 45152 38004
rect 40040 37884 40092 37936
rect 45100 37961 45109 37995
rect 45109 37961 45143 37995
rect 45143 37961 45152 37995
rect 45100 37952 45152 37961
rect 46112 37995 46164 38004
rect 46112 37961 46121 37995
rect 46121 37961 46155 37995
rect 46155 37961 46164 37995
rect 46112 37952 46164 37961
rect 46848 37995 46900 38004
rect 46848 37961 46857 37995
rect 46857 37961 46891 37995
rect 46891 37961 46900 37995
rect 46848 37952 46900 37961
rect 31024 37791 31076 37800
rect 31024 37757 31033 37791
rect 31033 37757 31067 37791
rect 31067 37757 31076 37791
rect 31024 37748 31076 37757
rect 37464 37791 37516 37800
rect 37464 37757 37473 37791
rect 37473 37757 37507 37791
rect 37507 37757 37516 37791
rect 37464 37748 37516 37757
rect 33968 37655 34020 37664
rect 33968 37621 33977 37655
rect 33977 37621 34011 37655
rect 34011 37621 34020 37655
rect 33968 37612 34020 37621
rect 37464 37612 37516 37664
rect 38108 37612 38160 37664
rect 44272 37816 44324 37868
rect 46296 37859 46348 37868
rect 46296 37825 46305 37859
rect 46305 37825 46339 37859
rect 46339 37825 46348 37859
rect 46296 37816 46348 37825
rect 46756 37859 46808 37868
rect 46756 37825 46765 37859
rect 46765 37825 46799 37859
rect 46799 37825 46808 37859
rect 46756 37816 46808 37825
rect 47308 37816 47360 37868
rect 47676 37816 47728 37868
rect 43076 37748 43128 37800
rect 43352 37748 43404 37800
rect 40316 37612 40368 37664
rect 41052 37655 41104 37664
rect 41052 37621 41061 37655
rect 41061 37621 41095 37655
rect 41095 37621 41104 37655
rect 41052 37612 41104 37621
rect 42892 37612 42944 37664
rect 47400 37612 47452 37664
rect 47860 37655 47912 37664
rect 47860 37621 47869 37655
rect 47869 37621 47903 37655
rect 47903 37621 47912 37655
rect 47860 37612 47912 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 24768 37408 24820 37460
rect 31024 37408 31076 37460
rect 35440 37408 35492 37460
rect 25320 37340 25372 37392
rect 26056 37340 26108 37392
rect 26240 37383 26292 37392
rect 26240 37349 26249 37383
rect 26249 37349 26283 37383
rect 26283 37349 26292 37383
rect 26240 37340 26292 37349
rect 33048 37383 33100 37392
rect 33048 37349 33057 37383
rect 33057 37349 33091 37383
rect 33091 37349 33100 37383
rect 33048 37340 33100 37349
rect 34612 37340 34664 37392
rect 24952 37272 25004 37324
rect 27528 37272 27580 37324
rect 27988 37315 28040 37324
rect 27988 37281 27997 37315
rect 27997 37281 28031 37315
rect 28031 37281 28040 37315
rect 27988 37272 28040 37281
rect 34704 37272 34756 37324
rect 35532 37315 35584 37324
rect 35532 37281 35541 37315
rect 35541 37281 35575 37315
rect 35575 37281 35584 37315
rect 35532 37272 35584 37281
rect 24676 37204 24728 37256
rect 26056 37247 26108 37256
rect 26056 37213 26065 37247
rect 26065 37213 26099 37247
rect 26099 37213 26108 37247
rect 26056 37204 26108 37213
rect 26332 37247 26384 37256
rect 26332 37213 26341 37247
rect 26341 37213 26375 37247
rect 26375 37213 26384 37247
rect 26332 37204 26384 37213
rect 28172 37247 28224 37256
rect 28172 37213 28181 37247
rect 28181 37213 28215 37247
rect 28215 37213 28224 37247
rect 28172 37204 28224 37213
rect 32128 37204 32180 37256
rect 32312 37247 32364 37256
rect 32312 37213 32321 37247
rect 32321 37213 32355 37247
rect 32355 37213 32364 37247
rect 32312 37204 32364 37213
rect 33324 37247 33376 37256
rect 33324 37213 33333 37247
rect 33333 37213 33367 37247
rect 33367 37213 33376 37247
rect 33324 37204 33376 37213
rect 33968 37204 34020 37256
rect 34796 37204 34848 37256
rect 37280 37408 37332 37460
rect 37924 37451 37976 37460
rect 37924 37417 37933 37451
rect 37933 37417 37967 37451
rect 37967 37417 37976 37451
rect 37924 37408 37976 37417
rect 42800 37408 42852 37460
rect 46296 37408 46348 37460
rect 41052 37272 41104 37324
rect 46204 37340 46256 37392
rect 44180 37272 44232 37324
rect 48228 37315 48280 37324
rect 48228 37281 48237 37315
rect 48237 37281 48271 37315
rect 48271 37281 48280 37315
rect 48228 37272 48280 37281
rect 36820 37204 36872 37256
rect 37188 37204 37240 37256
rect 40040 37247 40092 37256
rect 40040 37213 40049 37247
rect 40049 37213 40083 37247
rect 40083 37213 40092 37247
rect 40040 37204 40092 37213
rect 40316 37247 40368 37256
rect 40316 37213 40325 37247
rect 40325 37213 40359 37247
rect 40359 37213 40368 37247
rect 40316 37204 40368 37213
rect 26608 37136 26660 37188
rect 28908 37136 28960 37188
rect 23388 37068 23440 37120
rect 26240 37068 26292 37120
rect 28448 37068 28500 37120
rect 33140 37136 33192 37188
rect 33416 37179 33468 37188
rect 33416 37145 33425 37179
rect 33425 37145 33459 37179
rect 33459 37145 33468 37179
rect 33416 37136 33468 37145
rect 33232 37111 33284 37120
rect 33232 37077 33241 37111
rect 33241 37077 33275 37111
rect 33275 37077 33284 37111
rect 33232 37068 33284 37077
rect 34888 37111 34940 37120
rect 34888 37077 34897 37111
rect 34897 37077 34931 37111
rect 34931 37077 34940 37111
rect 34888 37068 34940 37077
rect 35256 37179 35308 37188
rect 35256 37145 35265 37179
rect 35265 37145 35299 37179
rect 35299 37145 35308 37179
rect 35256 37136 35308 37145
rect 36176 37136 36228 37188
rect 37556 37136 37608 37188
rect 39948 37136 40000 37188
rect 35900 37068 35952 37120
rect 36452 37068 36504 37120
rect 40960 37068 41012 37120
rect 43352 37204 43404 37256
rect 44088 37247 44140 37256
rect 44088 37213 44097 37247
rect 44097 37213 44131 37247
rect 44131 37213 44140 37247
rect 44088 37204 44140 37213
rect 44272 37247 44324 37256
rect 44272 37213 44281 37247
rect 44281 37213 44315 37247
rect 44315 37213 44324 37247
rect 44272 37204 44324 37213
rect 41420 37179 41472 37188
rect 41420 37145 41429 37179
rect 41429 37145 41463 37179
rect 41463 37145 41472 37179
rect 41420 37136 41472 37145
rect 42616 37136 42668 37188
rect 45376 37136 45428 37188
rect 45836 37068 45888 37120
rect 47860 37136 47912 37188
rect 47952 37068 48004 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 25964 36864 26016 36916
rect 28172 36864 28224 36916
rect 24952 36839 25004 36848
rect 24952 36805 24961 36839
rect 24961 36805 24995 36839
rect 24995 36805 25004 36839
rect 24952 36796 25004 36805
rect 25780 36796 25832 36848
rect 26148 36839 26200 36848
rect 26148 36805 26157 36839
rect 26157 36805 26191 36839
rect 26191 36805 26200 36839
rect 26148 36796 26200 36805
rect 26240 36839 26292 36848
rect 26240 36805 26275 36839
rect 26275 36805 26292 36839
rect 26240 36796 26292 36805
rect 26976 36796 27028 36848
rect 32312 36864 32364 36916
rect 36176 36907 36228 36916
rect 24676 36728 24728 36780
rect 24032 36524 24084 36576
rect 28264 36728 28316 36780
rect 26608 36660 26660 36712
rect 27160 36703 27212 36712
rect 27160 36669 27169 36703
rect 27169 36669 27203 36703
rect 27203 36669 27212 36703
rect 27160 36660 27212 36669
rect 26056 36592 26108 36644
rect 25780 36567 25832 36576
rect 25780 36533 25789 36567
rect 25789 36533 25823 36567
rect 25823 36533 25832 36567
rect 25780 36524 25832 36533
rect 25872 36524 25924 36576
rect 27344 36524 27396 36576
rect 32036 36796 32088 36848
rect 32128 36796 32180 36848
rect 30656 36728 30708 36780
rect 31208 36728 31260 36780
rect 33140 36771 33192 36780
rect 33140 36737 33149 36771
rect 33149 36737 33183 36771
rect 33183 36737 33192 36771
rect 33140 36728 33192 36737
rect 33324 36771 33376 36780
rect 33324 36737 33333 36771
rect 33333 36737 33367 36771
rect 33367 36737 33376 36771
rect 33324 36728 33376 36737
rect 34888 36796 34940 36848
rect 35624 36796 35676 36848
rect 36176 36873 36185 36907
rect 36185 36873 36219 36907
rect 36219 36873 36228 36907
rect 36176 36864 36228 36873
rect 37464 36864 37516 36916
rect 42616 36907 42668 36916
rect 42616 36873 42625 36907
rect 42625 36873 42659 36907
rect 42659 36873 42668 36907
rect 42616 36864 42668 36873
rect 33048 36660 33100 36712
rect 35348 36728 35400 36780
rect 36452 36771 36504 36780
rect 36452 36737 36461 36771
rect 36461 36737 36495 36771
rect 36495 36737 36504 36771
rect 36728 36796 36780 36848
rect 39028 36839 39080 36848
rect 39028 36805 39037 36839
rect 39037 36805 39071 36839
rect 39071 36805 39080 36839
rect 39028 36796 39080 36805
rect 39212 36796 39264 36848
rect 47676 36796 47728 36848
rect 36452 36728 36504 36737
rect 37556 36728 37608 36780
rect 41052 36728 41104 36780
rect 42800 36771 42852 36780
rect 42800 36737 42809 36771
rect 42809 36737 42843 36771
rect 42843 36737 42852 36771
rect 42800 36728 42852 36737
rect 37280 36660 37332 36712
rect 38568 36660 38620 36712
rect 40316 36660 40368 36712
rect 41144 36660 41196 36712
rect 33140 36524 33192 36576
rect 33232 36524 33284 36576
rect 33416 36567 33468 36576
rect 33416 36533 33425 36567
rect 33425 36533 33459 36567
rect 33459 36533 33468 36567
rect 33416 36524 33468 36533
rect 37832 36567 37884 36576
rect 37832 36533 37841 36567
rect 37841 36533 37875 36567
rect 37875 36533 37884 36567
rect 37832 36524 37884 36533
rect 39672 36524 39724 36576
rect 46480 36524 46532 36576
rect 47860 36567 47912 36576
rect 47860 36533 47869 36567
rect 47869 36533 47903 36567
rect 47903 36533 47912 36567
rect 47860 36524 47912 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 28264 36363 28316 36372
rect 28264 36329 28273 36363
rect 28273 36329 28307 36363
rect 28307 36329 28316 36363
rect 28264 36320 28316 36329
rect 32128 36320 32180 36372
rect 33140 36320 33192 36372
rect 39212 36320 39264 36372
rect 39948 36252 40000 36304
rect 40040 36252 40092 36304
rect 37188 36184 37240 36236
rect 39028 36184 39080 36236
rect 46480 36227 46532 36236
rect 23388 36159 23440 36168
rect 23388 36125 23397 36159
rect 23397 36125 23431 36159
rect 23431 36125 23440 36159
rect 23388 36116 23440 36125
rect 24032 36159 24084 36168
rect 24032 36125 24041 36159
rect 24041 36125 24075 36159
rect 24075 36125 24084 36159
rect 24032 36116 24084 36125
rect 28448 36159 28500 36168
rect 28448 36125 28457 36159
rect 28457 36125 28491 36159
rect 28491 36125 28500 36159
rect 28448 36116 28500 36125
rect 34520 36116 34572 36168
rect 37464 36116 37516 36168
rect 39948 36116 40000 36168
rect 41052 36116 41104 36168
rect 41144 36159 41196 36168
rect 41144 36125 41153 36159
rect 41153 36125 41187 36159
rect 41187 36125 41196 36159
rect 46480 36193 46489 36227
rect 46489 36193 46523 36227
rect 46523 36193 46532 36227
rect 46480 36184 46532 36193
rect 47860 36184 47912 36236
rect 48228 36227 48280 36236
rect 48228 36193 48237 36227
rect 48237 36193 48271 36227
rect 48271 36193 48280 36227
rect 48228 36184 48280 36193
rect 41144 36116 41196 36125
rect 44180 36116 44232 36168
rect 23756 35980 23808 36032
rect 24032 35980 24084 36032
rect 26240 35980 26292 36032
rect 27160 35980 27212 36032
rect 35900 36048 35952 36100
rect 43352 36091 43404 36100
rect 43352 36057 43361 36091
rect 43361 36057 43395 36091
rect 43395 36057 43404 36091
rect 43352 36048 43404 36057
rect 43996 36048 44048 36100
rect 36728 35980 36780 36032
rect 36820 36023 36872 36032
rect 36820 35989 36829 36023
rect 36829 35989 36863 36023
rect 36863 35989 36872 36023
rect 36820 35980 36872 35989
rect 39580 35980 39632 36032
rect 40500 36023 40552 36032
rect 40500 35989 40509 36023
rect 40509 35989 40543 36023
rect 40543 35989 40552 36023
rect 40500 35980 40552 35989
rect 40684 35980 40736 36032
rect 44180 36023 44232 36032
rect 44180 35989 44189 36023
rect 44189 35989 44223 36023
rect 44223 35989 44232 36023
rect 44180 35980 44232 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 25964 35819 26016 35828
rect 25964 35785 25973 35819
rect 25973 35785 26007 35819
rect 26007 35785 26016 35819
rect 25964 35776 26016 35785
rect 27528 35819 27580 35828
rect 27528 35785 27537 35819
rect 27537 35785 27571 35819
rect 27571 35785 27580 35819
rect 27528 35776 27580 35785
rect 33416 35776 33468 35828
rect 34704 35819 34756 35828
rect 34704 35785 34729 35819
rect 34729 35785 34756 35819
rect 34888 35819 34940 35828
rect 34704 35776 34756 35785
rect 34888 35785 34897 35819
rect 34897 35785 34931 35819
rect 34931 35785 34940 35819
rect 34888 35776 34940 35785
rect 35900 35819 35952 35828
rect 35900 35785 35909 35819
rect 35909 35785 35943 35819
rect 35943 35785 35952 35819
rect 35900 35776 35952 35785
rect 23756 35708 23808 35760
rect 25320 35640 25372 35692
rect 27344 35683 27396 35692
rect 27344 35649 27353 35683
rect 27353 35649 27387 35683
rect 27387 35649 27396 35683
rect 27344 35640 27396 35649
rect 28080 35640 28132 35692
rect 29276 35640 29328 35692
rect 32128 35640 32180 35692
rect 32588 35683 32640 35692
rect 32588 35649 32622 35683
rect 32622 35649 32640 35683
rect 32588 35640 32640 35649
rect 33692 35640 33744 35692
rect 36820 35708 36872 35760
rect 37832 35640 37884 35692
rect 39488 35776 39540 35828
rect 40684 35776 40736 35828
rect 41328 35776 41380 35828
rect 42800 35776 42852 35828
rect 43260 35776 43312 35828
rect 39304 35683 39356 35692
rect 24584 35615 24636 35624
rect 24584 35581 24593 35615
rect 24593 35581 24627 35615
rect 24627 35581 24636 35615
rect 24584 35572 24636 35581
rect 39304 35649 39313 35683
rect 39313 35649 39347 35683
rect 39347 35649 39356 35683
rect 39304 35640 39356 35649
rect 39488 35683 39540 35692
rect 39488 35649 39497 35683
rect 39497 35649 39531 35683
rect 39531 35649 39540 35683
rect 39488 35640 39540 35649
rect 39580 35683 39632 35692
rect 39580 35649 39589 35683
rect 39589 35649 39623 35683
rect 39623 35649 39632 35683
rect 40500 35708 40552 35760
rect 39580 35640 39632 35649
rect 40684 35683 40736 35692
rect 40684 35649 40693 35683
rect 40693 35649 40727 35683
rect 40727 35649 40736 35683
rect 40684 35640 40736 35649
rect 40960 35683 41012 35692
rect 40960 35649 40969 35683
rect 40969 35649 41003 35683
rect 41003 35649 41012 35683
rect 40960 35640 41012 35649
rect 41052 35683 41104 35692
rect 41052 35649 41061 35683
rect 41061 35649 41095 35683
rect 41095 35649 41104 35683
rect 43352 35708 43404 35760
rect 44272 35776 44324 35828
rect 47124 35708 47176 35760
rect 41052 35640 41104 35649
rect 39672 35615 39724 35624
rect 39672 35581 39681 35615
rect 39681 35581 39715 35615
rect 39715 35581 39724 35615
rect 39672 35572 39724 35581
rect 27988 35436 28040 35488
rect 30564 35479 30616 35488
rect 30564 35445 30573 35479
rect 30573 35445 30607 35479
rect 30607 35445 30616 35479
rect 30564 35436 30616 35445
rect 34796 35436 34848 35488
rect 35348 35436 35400 35488
rect 38568 35436 38620 35488
rect 39304 35436 39356 35488
rect 41052 35504 41104 35556
rect 40040 35479 40092 35488
rect 40040 35445 40049 35479
rect 40049 35445 40083 35479
rect 40083 35445 40092 35479
rect 40040 35436 40092 35445
rect 40500 35479 40552 35488
rect 40500 35445 40509 35479
rect 40509 35445 40543 35479
rect 40543 35445 40552 35479
rect 40500 35436 40552 35445
rect 42892 35640 42944 35692
rect 45192 35640 45244 35692
rect 46664 35683 46716 35692
rect 46664 35649 46673 35683
rect 46673 35649 46707 35683
rect 46707 35649 46716 35683
rect 46664 35640 46716 35649
rect 47216 35640 47268 35692
rect 44364 35572 44416 35624
rect 48136 35504 48188 35556
rect 44364 35436 44416 35488
rect 47032 35436 47084 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 26332 35232 26384 35284
rect 26700 35232 26752 35284
rect 29276 35232 29328 35284
rect 32588 35232 32640 35284
rect 42892 35275 42944 35284
rect 42892 35241 42901 35275
rect 42901 35241 42935 35275
rect 42935 35241 42944 35275
rect 42892 35232 42944 35241
rect 24584 35028 24636 35080
rect 30564 35139 30616 35148
rect 30564 35105 30573 35139
rect 30573 35105 30607 35139
rect 30607 35105 30616 35139
rect 30564 35096 30616 35105
rect 25780 34960 25832 35012
rect 30472 35028 30524 35080
rect 33232 35071 33284 35080
rect 30380 34960 30432 35012
rect 33232 35037 33241 35071
rect 33241 35037 33275 35071
rect 33275 35037 33284 35071
rect 33232 35028 33284 35037
rect 38568 35071 38620 35080
rect 38568 35037 38577 35071
rect 38577 35037 38611 35071
rect 38611 35037 38620 35071
rect 38568 35028 38620 35037
rect 40960 35096 41012 35148
rect 40408 35071 40460 35080
rect 40408 35037 40417 35071
rect 40417 35037 40451 35071
rect 40451 35037 40460 35071
rect 40408 35028 40460 35037
rect 40684 35028 40736 35080
rect 43168 35071 43220 35080
rect 43168 35037 43177 35071
rect 43177 35037 43211 35071
rect 43211 35037 43220 35071
rect 43168 35028 43220 35037
rect 43352 35164 43404 35216
rect 44548 35096 44600 35148
rect 45192 35096 45244 35148
rect 45928 35139 45980 35148
rect 45928 35105 45937 35139
rect 45937 35105 45971 35139
rect 45971 35105 45980 35139
rect 45928 35096 45980 35105
rect 43444 35028 43496 35080
rect 43536 35071 43588 35080
rect 43536 35037 43545 35071
rect 43545 35037 43579 35071
rect 43579 35037 43588 35071
rect 44180 35071 44232 35080
rect 43536 35028 43588 35037
rect 44180 35037 44189 35071
rect 44189 35037 44223 35071
rect 44223 35037 44232 35071
rect 44180 35028 44232 35037
rect 46020 35028 46072 35080
rect 46940 35071 46992 35080
rect 46940 35037 46949 35071
rect 46949 35037 46983 35071
rect 46983 35037 46992 35071
rect 46940 35028 46992 35037
rect 47032 35028 47084 35080
rect 33876 34960 33928 35012
rect 39120 34960 39172 35012
rect 42800 34960 42852 35012
rect 26056 34892 26108 34944
rect 31392 34935 31444 34944
rect 31392 34901 31401 34935
rect 31401 34901 31435 34935
rect 31435 34901 31444 34935
rect 31392 34892 31444 34901
rect 38016 34935 38068 34944
rect 38016 34901 38025 34935
rect 38025 34901 38059 34935
rect 38059 34901 38068 34935
rect 38016 34892 38068 34901
rect 40132 34892 40184 34944
rect 46848 34892 46900 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 25320 34731 25372 34740
rect 25320 34697 25329 34731
rect 25329 34697 25363 34731
rect 25363 34697 25372 34731
rect 25320 34688 25372 34697
rect 30380 34688 30432 34740
rect 31116 34688 31168 34740
rect 33232 34688 33284 34740
rect 35440 34688 35492 34740
rect 24584 34620 24636 34672
rect 24032 34552 24084 34604
rect 27528 34620 27580 34672
rect 29460 34620 29512 34672
rect 27436 34552 27488 34604
rect 28080 34552 28132 34604
rect 28908 34552 28960 34604
rect 32128 34620 32180 34672
rect 43444 34688 43496 34740
rect 44180 34688 44232 34740
rect 46664 34688 46716 34740
rect 31392 34552 31444 34604
rect 33692 34595 33744 34604
rect 33692 34561 33701 34595
rect 33701 34561 33735 34595
rect 33735 34561 33744 34595
rect 33692 34552 33744 34561
rect 33876 34595 33928 34604
rect 33876 34561 33885 34595
rect 33885 34561 33919 34595
rect 33919 34561 33928 34595
rect 33876 34552 33928 34561
rect 34520 34595 34572 34604
rect 34520 34561 34529 34595
rect 34529 34561 34563 34595
rect 34563 34561 34572 34595
rect 34520 34552 34572 34561
rect 35716 34552 35768 34604
rect 38292 34552 38344 34604
rect 38752 34552 38804 34604
rect 40040 34620 40092 34672
rect 40132 34620 40184 34672
rect 40500 34552 40552 34604
rect 38936 34484 38988 34536
rect 39396 34484 39448 34536
rect 43260 34552 43312 34604
rect 44272 34595 44324 34604
rect 44272 34561 44281 34595
rect 44281 34561 44315 34595
rect 44315 34561 44324 34595
rect 44272 34552 44324 34561
rect 44548 34595 44600 34604
rect 44548 34561 44557 34595
rect 44557 34561 44591 34595
rect 44591 34561 44600 34595
rect 44548 34552 44600 34561
rect 46020 34552 46072 34604
rect 46848 34595 46900 34604
rect 46848 34561 46857 34595
rect 46857 34561 46891 34595
rect 46891 34561 46900 34595
rect 46848 34552 46900 34561
rect 38016 34416 38068 34468
rect 38844 34416 38896 34468
rect 44180 34484 44232 34536
rect 44364 34484 44416 34536
rect 45928 34527 45980 34536
rect 45928 34493 45937 34527
rect 45937 34493 45971 34527
rect 45971 34493 45980 34527
rect 45928 34484 45980 34493
rect 47400 34484 47452 34536
rect 27344 34348 27396 34400
rect 31760 34391 31812 34400
rect 31760 34357 31769 34391
rect 31769 34357 31803 34391
rect 31803 34357 31812 34391
rect 31760 34348 31812 34357
rect 34336 34348 34388 34400
rect 37096 34348 37148 34400
rect 41328 34416 41380 34468
rect 47216 34416 47268 34468
rect 40684 34348 40736 34400
rect 47124 34348 47176 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 28908 34187 28960 34196
rect 28908 34153 28917 34187
rect 28917 34153 28951 34187
rect 28951 34153 28960 34187
rect 28908 34144 28960 34153
rect 35716 34187 35768 34196
rect 35716 34153 35725 34187
rect 35725 34153 35759 34187
rect 35759 34153 35768 34187
rect 35716 34144 35768 34153
rect 43996 34187 44048 34196
rect 43996 34153 44005 34187
rect 44005 34153 44039 34187
rect 44039 34153 44048 34187
rect 43996 34144 44048 34153
rect 48136 34187 48188 34196
rect 48136 34153 48145 34187
rect 48145 34153 48179 34187
rect 48179 34153 48188 34187
rect 48136 34144 48188 34153
rect 33876 34076 33928 34128
rect 26056 33983 26108 33992
rect 26056 33949 26065 33983
rect 26065 33949 26099 33983
rect 26099 33949 26108 33983
rect 26056 33940 26108 33949
rect 34520 34008 34572 34060
rect 37740 34008 37792 34060
rect 38292 34076 38344 34128
rect 29828 33983 29880 33992
rect 29828 33949 29837 33983
rect 29837 33949 29871 33983
rect 29871 33949 29880 33983
rect 29828 33940 29880 33949
rect 30380 33940 30432 33992
rect 30564 33940 30616 33992
rect 27160 33872 27212 33924
rect 31760 33940 31812 33992
rect 34336 33983 34388 33992
rect 34336 33949 34345 33983
rect 34345 33949 34379 33983
rect 34379 33949 34388 33983
rect 34336 33940 34388 33949
rect 34796 33940 34848 33992
rect 38936 33983 38988 33992
rect 33508 33915 33560 33924
rect 33508 33881 33517 33915
rect 33517 33881 33551 33915
rect 33551 33881 33560 33915
rect 33508 33872 33560 33881
rect 33876 33872 33928 33924
rect 37464 33872 37516 33924
rect 38936 33949 38945 33983
rect 38945 33949 38979 33983
rect 38979 33949 38988 33983
rect 38936 33940 38988 33949
rect 39028 33983 39080 33992
rect 39028 33949 39037 33983
rect 39037 33949 39071 33983
rect 39071 33949 39080 33983
rect 39028 33940 39080 33949
rect 39120 33872 39172 33924
rect 40040 33983 40092 33992
rect 40040 33949 40049 33983
rect 40049 33949 40083 33983
rect 40083 33949 40092 33983
rect 40040 33940 40092 33949
rect 40684 33983 40736 33992
rect 40684 33949 40693 33983
rect 40693 33949 40727 33983
rect 40727 33949 40736 33983
rect 40684 33940 40736 33949
rect 40500 33872 40552 33924
rect 41052 33940 41104 33992
rect 44180 33983 44232 33992
rect 44180 33949 44189 33983
rect 44189 33949 44223 33983
rect 44223 33949 44232 33983
rect 44180 33940 44232 33949
rect 45376 33940 45428 33992
rect 48320 33983 48372 33992
rect 48320 33949 48329 33983
rect 48329 33949 48363 33983
rect 48363 33949 48372 33983
rect 48320 33940 48372 33949
rect 27068 33804 27120 33856
rect 31116 33847 31168 33856
rect 31116 33813 31125 33847
rect 31125 33813 31159 33847
rect 31159 33813 31168 33847
rect 31116 33804 31168 33813
rect 32496 33804 32548 33856
rect 34520 33804 34572 33856
rect 38200 33804 38252 33856
rect 44180 33804 44232 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 27160 33643 27212 33652
rect 27160 33609 27169 33643
rect 27169 33609 27203 33643
rect 27203 33609 27212 33643
rect 27160 33600 27212 33609
rect 24952 33464 25004 33516
rect 27436 33532 27488 33584
rect 30564 33532 30616 33584
rect 32128 33532 32180 33584
rect 34520 33575 34572 33584
rect 27344 33507 27396 33516
rect 27344 33473 27353 33507
rect 27353 33473 27387 33507
rect 27387 33473 27396 33507
rect 27344 33464 27396 33473
rect 29828 33464 29880 33516
rect 33508 33464 33560 33516
rect 34520 33541 34554 33575
rect 34554 33541 34572 33575
rect 34520 33532 34572 33541
rect 34796 33600 34848 33652
rect 37464 33643 37516 33652
rect 37464 33609 37473 33643
rect 37473 33609 37507 33643
rect 37507 33609 37516 33643
rect 37464 33600 37516 33609
rect 37096 33532 37148 33584
rect 26700 33396 26752 33448
rect 31760 33396 31812 33448
rect 33416 33439 33468 33448
rect 33416 33405 33425 33439
rect 33425 33405 33459 33439
rect 33459 33405 33468 33439
rect 33416 33396 33468 33405
rect 37556 33464 37608 33516
rect 37740 33507 37792 33516
rect 37740 33473 37749 33507
rect 37749 33473 37783 33507
rect 37783 33473 37792 33507
rect 37740 33464 37792 33473
rect 38016 33600 38068 33652
rect 39028 33600 39080 33652
rect 38200 33532 38252 33584
rect 38292 33464 38344 33516
rect 38752 33507 38804 33516
rect 38752 33473 38761 33507
rect 38761 33473 38795 33507
rect 38795 33473 38804 33507
rect 38752 33464 38804 33473
rect 38936 33396 38988 33448
rect 41420 33600 41472 33652
rect 41236 33532 41288 33584
rect 40868 33464 40920 33516
rect 45100 33464 45152 33516
rect 44180 33396 44232 33448
rect 45192 33439 45244 33448
rect 45192 33405 45201 33439
rect 45201 33405 45235 33439
rect 45235 33405 45244 33439
rect 45192 33396 45244 33405
rect 41052 33328 41104 33380
rect 2320 33303 2372 33312
rect 2320 33269 2329 33303
rect 2329 33269 2363 33303
rect 2363 33269 2372 33303
rect 2320 33260 2372 33269
rect 24860 33260 24912 33312
rect 31116 33303 31168 33312
rect 31116 33269 31125 33303
rect 31125 33269 31159 33303
rect 31159 33269 31168 33303
rect 31116 33260 31168 33269
rect 31392 33303 31444 33312
rect 31392 33269 31401 33303
rect 31401 33269 31435 33303
rect 31435 33269 31444 33303
rect 31392 33260 31444 33269
rect 34152 33260 34204 33312
rect 41144 33260 41196 33312
rect 45284 33260 45336 33312
rect 47952 33303 48004 33312
rect 47952 33269 47961 33303
rect 47961 33269 47995 33303
rect 47995 33269 48004 33303
rect 47952 33260 48004 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 39120 33056 39172 33108
rect 43168 33056 43220 33108
rect 44548 33056 44600 33108
rect 25964 32988 26016 33040
rect 26700 33031 26752 33040
rect 26700 32997 26709 33031
rect 26709 32997 26743 33031
rect 26743 32997 26752 33031
rect 26700 32988 26752 32997
rect 2320 32920 2372 32972
rect 2780 32963 2832 32972
rect 2780 32929 2789 32963
rect 2789 32929 2823 32963
rect 2823 32929 2832 32963
rect 2780 32920 2832 32929
rect 32128 32963 32180 32972
rect 32128 32929 32137 32963
rect 32137 32929 32171 32963
rect 32171 32929 32180 32963
rect 32128 32920 32180 32929
rect 26056 32852 26108 32904
rect 30564 32852 30616 32904
rect 31392 32852 31444 32904
rect 34152 32895 34204 32904
rect 34152 32861 34161 32895
rect 34161 32861 34195 32895
rect 34195 32861 34204 32895
rect 34152 32852 34204 32861
rect 40040 32920 40092 32972
rect 41052 32920 41104 32972
rect 42616 32920 42668 32972
rect 44180 32988 44232 33040
rect 43904 32963 43956 32972
rect 43904 32929 43913 32963
rect 43913 32929 43947 32963
rect 43947 32929 43956 32963
rect 43904 32920 43956 32929
rect 2412 32784 2464 32836
rect 24860 32827 24912 32836
rect 24860 32793 24894 32827
rect 24894 32793 24912 32827
rect 24860 32784 24912 32793
rect 26424 32827 26476 32836
rect 26424 32793 26433 32827
rect 26433 32793 26467 32827
rect 26467 32793 26476 32827
rect 26424 32784 26476 32793
rect 27528 32784 27580 32836
rect 31760 32784 31812 32836
rect 32404 32827 32456 32836
rect 32404 32793 32438 32827
rect 32438 32793 32456 32827
rect 32404 32784 32456 32793
rect 37188 32784 37240 32836
rect 37280 32784 37332 32836
rect 40868 32784 40920 32836
rect 43352 32852 43404 32904
rect 43536 32895 43588 32904
rect 43536 32861 43545 32895
rect 43545 32861 43579 32895
rect 43579 32861 43588 32895
rect 43536 32852 43588 32861
rect 45284 32920 45336 32972
rect 47952 32920 48004 32972
rect 44548 32895 44600 32904
rect 44548 32861 44557 32895
rect 44557 32861 44591 32895
rect 44591 32861 44600 32895
rect 44548 32852 44600 32861
rect 45652 32895 45704 32904
rect 45652 32861 45661 32895
rect 45661 32861 45695 32895
rect 45695 32861 45704 32895
rect 45652 32852 45704 32861
rect 41788 32827 41840 32836
rect 41788 32793 41822 32827
rect 41822 32793 41840 32827
rect 41788 32784 41840 32793
rect 47860 32784 47912 32836
rect 48320 32827 48372 32836
rect 48320 32793 48329 32827
rect 48329 32793 48363 32827
rect 48363 32793 48372 32827
rect 48320 32784 48372 32793
rect 26240 32716 26292 32768
rect 26884 32759 26936 32768
rect 26884 32725 26893 32759
rect 26893 32725 26927 32759
rect 26927 32725 26936 32759
rect 26884 32716 26936 32725
rect 29736 32759 29788 32768
rect 29736 32725 29745 32759
rect 29745 32725 29779 32759
rect 29779 32725 29788 32759
rect 29736 32716 29788 32725
rect 32772 32716 32824 32768
rect 33416 32716 33468 32768
rect 33968 32759 34020 32768
rect 33968 32725 33977 32759
rect 33977 32725 34011 32759
rect 34011 32725 34020 32759
rect 33968 32716 34020 32725
rect 37740 32759 37792 32768
rect 37740 32725 37749 32759
rect 37749 32725 37783 32759
rect 37783 32725 37792 32759
rect 37740 32716 37792 32725
rect 38660 32716 38712 32768
rect 40316 32716 40368 32768
rect 41328 32716 41380 32768
rect 44824 32716 44876 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 2412 32555 2464 32564
rect 2412 32521 2421 32555
rect 2421 32521 2455 32555
rect 2455 32521 2464 32555
rect 2412 32512 2464 32521
rect 10508 32444 10560 32496
rect 2596 32376 2648 32428
rect 7380 32376 7432 32428
rect 27068 32512 27120 32564
rect 29828 32512 29880 32564
rect 32404 32512 32456 32564
rect 32496 32512 32548 32564
rect 25964 32419 26016 32428
rect 25964 32385 25973 32419
rect 25973 32385 26007 32419
rect 26007 32385 26016 32419
rect 25964 32376 26016 32385
rect 26056 32376 26108 32428
rect 29736 32444 29788 32496
rect 32772 32487 32824 32496
rect 32772 32453 32807 32487
rect 32807 32453 32824 32487
rect 32772 32444 32824 32453
rect 26240 32351 26292 32360
rect 26240 32317 26249 32351
rect 26249 32317 26283 32351
rect 26283 32317 26292 32351
rect 26240 32308 26292 32317
rect 26424 32351 26476 32360
rect 26424 32317 26458 32351
rect 26458 32317 26476 32351
rect 26424 32308 26476 32317
rect 26700 32308 26752 32360
rect 27252 32240 27304 32292
rect 27528 32283 27580 32292
rect 27528 32249 27537 32283
rect 27537 32249 27571 32283
rect 27571 32249 27580 32283
rect 27528 32240 27580 32249
rect 32404 32376 32456 32428
rect 33968 32376 34020 32428
rect 32772 32308 32824 32360
rect 35532 32308 35584 32360
rect 41604 32512 41656 32564
rect 41788 32512 41840 32564
rect 41880 32512 41932 32564
rect 43260 32512 43312 32564
rect 44824 32555 44876 32564
rect 44824 32521 44833 32555
rect 44833 32521 44867 32555
rect 44867 32521 44876 32555
rect 44824 32512 44876 32521
rect 45284 32512 45336 32564
rect 47860 32555 47912 32564
rect 37464 32419 37516 32428
rect 37464 32385 37473 32419
rect 37473 32385 37507 32419
rect 37507 32385 37516 32419
rect 37464 32376 37516 32385
rect 37556 32376 37608 32428
rect 39120 32444 39172 32496
rect 39212 32376 39264 32428
rect 40040 32376 40092 32428
rect 41052 32444 41104 32496
rect 41236 32444 41288 32496
rect 37188 32240 37240 32292
rect 40040 32240 40092 32292
rect 40408 32351 40460 32360
rect 40408 32317 40417 32351
rect 40417 32317 40451 32351
rect 40451 32317 40460 32351
rect 40408 32308 40460 32317
rect 40592 32240 40644 32292
rect 41144 32419 41196 32428
rect 41144 32385 41153 32419
rect 41153 32385 41187 32419
rect 41187 32385 41196 32419
rect 41144 32376 41196 32385
rect 41420 32376 41472 32428
rect 41696 32376 41748 32428
rect 42616 32419 42668 32428
rect 42616 32385 42625 32419
rect 42625 32385 42659 32419
rect 42659 32385 42668 32419
rect 42616 32376 42668 32385
rect 40868 32308 40920 32360
rect 41880 32308 41932 32360
rect 42708 32240 42760 32292
rect 26240 32172 26292 32224
rect 26792 32172 26844 32224
rect 27620 32215 27672 32224
rect 27620 32181 27629 32215
rect 27629 32181 27663 32215
rect 27663 32181 27672 32215
rect 27620 32172 27672 32181
rect 40960 32172 41012 32224
rect 41144 32172 41196 32224
rect 43168 32376 43220 32428
rect 43812 32419 43864 32428
rect 43812 32385 43821 32419
rect 43821 32385 43855 32419
rect 43855 32385 43864 32419
rect 43812 32376 43864 32385
rect 45192 32444 45244 32496
rect 47860 32521 47869 32555
rect 47869 32521 47903 32555
rect 47903 32521 47912 32555
rect 47860 32512 47912 32521
rect 46664 32376 46716 32428
rect 47124 32376 47176 32428
rect 47860 32376 47912 32428
rect 48136 32376 48188 32428
rect 43536 32308 43588 32360
rect 44088 32308 44140 32360
rect 47400 32308 47452 32360
rect 46480 32283 46532 32292
rect 46480 32249 46489 32283
rect 46489 32249 46523 32283
rect 46523 32249 46532 32283
rect 46480 32240 46532 32249
rect 43352 32172 43404 32224
rect 47124 32215 47176 32224
rect 47124 32181 47133 32215
rect 47133 32181 47167 32215
rect 47167 32181 47176 32215
rect 47124 32172 47176 32181
rect 47400 32172 47452 32224
rect 47676 32172 47728 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 30564 32011 30616 32020
rect 30564 31977 30573 32011
rect 30573 31977 30607 32011
rect 30607 31977 30616 32011
rect 30564 31968 30616 31977
rect 36728 31968 36780 32020
rect 37188 31968 37240 32020
rect 37464 31968 37516 32020
rect 26332 31900 26384 31952
rect 26516 31764 26568 31816
rect 27068 31807 27120 31816
rect 27068 31773 27077 31807
rect 27077 31773 27111 31807
rect 27111 31773 27120 31807
rect 27068 31764 27120 31773
rect 27252 31807 27304 31816
rect 27252 31773 27261 31807
rect 27261 31773 27295 31807
rect 27295 31773 27304 31807
rect 27252 31764 27304 31773
rect 29092 31764 29144 31816
rect 30196 31807 30248 31816
rect 30196 31773 30205 31807
rect 30205 31773 30239 31807
rect 30239 31773 30248 31807
rect 30196 31764 30248 31773
rect 30380 31807 30432 31816
rect 30380 31773 30389 31807
rect 30389 31773 30423 31807
rect 30423 31773 30432 31807
rect 30380 31764 30432 31773
rect 37096 31900 37148 31952
rect 35624 31832 35676 31884
rect 37464 31832 37516 31884
rect 37740 31832 37792 31884
rect 38752 31900 38804 31952
rect 40316 31968 40368 32020
rect 40868 32011 40920 32020
rect 40868 31977 40877 32011
rect 40877 31977 40911 32011
rect 40911 31977 40920 32011
rect 40868 31968 40920 31977
rect 43812 31968 43864 32020
rect 45652 31968 45704 32020
rect 46664 31968 46716 32020
rect 40776 31900 40828 31952
rect 41052 31875 41104 31884
rect 35900 31764 35952 31816
rect 36084 31807 36136 31816
rect 36084 31773 36093 31807
rect 36093 31773 36127 31807
rect 36127 31773 36136 31807
rect 36084 31764 36136 31773
rect 38384 31764 38436 31816
rect 26792 31696 26844 31748
rect 26976 31696 27028 31748
rect 38568 31696 38620 31748
rect 38844 31764 38896 31816
rect 41052 31841 41061 31875
rect 41061 31841 41095 31875
rect 41095 31841 41104 31875
rect 41052 31832 41104 31841
rect 41236 31875 41288 31884
rect 41236 31841 41245 31875
rect 41245 31841 41279 31875
rect 41279 31841 41288 31875
rect 41236 31832 41288 31841
rect 43168 31900 43220 31952
rect 44088 31900 44140 31952
rect 45100 31832 45152 31884
rect 46664 31832 46716 31884
rect 46940 31875 46992 31884
rect 46940 31841 46949 31875
rect 46949 31841 46983 31875
rect 46983 31841 46992 31875
rect 46940 31832 46992 31841
rect 39396 31764 39448 31816
rect 40040 31807 40092 31816
rect 40040 31773 40049 31807
rect 40049 31773 40083 31807
rect 40083 31773 40092 31807
rect 40040 31764 40092 31773
rect 40592 31764 40644 31816
rect 40776 31764 40828 31816
rect 43904 31807 43956 31816
rect 43904 31773 43913 31807
rect 43913 31773 43947 31807
rect 43947 31773 43956 31807
rect 43904 31764 43956 31773
rect 45192 31764 45244 31816
rect 40960 31696 41012 31748
rect 44548 31696 44600 31748
rect 46940 31696 46992 31748
rect 26608 31628 26660 31680
rect 26884 31628 26936 31680
rect 27528 31628 27580 31680
rect 29736 31628 29788 31680
rect 39212 31628 39264 31680
rect 40592 31628 40644 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 26976 31424 27028 31476
rect 24952 31356 25004 31408
rect 24308 31288 24360 31340
rect 26240 31331 26292 31340
rect 26240 31297 26249 31331
rect 26249 31297 26283 31331
rect 26283 31297 26292 31331
rect 26240 31288 26292 31297
rect 26516 31288 26568 31340
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 27528 31356 27580 31408
rect 29736 31424 29788 31476
rect 26056 31127 26108 31136
rect 26056 31093 26065 31127
rect 26065 31093 26099 31127
rect 26099 31093 26108 31127
rect 26056 31084 26108 31093
rect 26608 31263 26660 31272
rect 26608 31229 26617 31263
rect 26617 31229 26651 31263
rect 26651 31229 26660 31263
rect 26608 31220 26660 31229
rect 27620 31288 27672 31340
rect 30196 31356 30248 31408
rect 30104 31288 30156 31340
rect 29092 31220 29144 31272
rect 29368 31263 29420 31272
rect 29368 31229 29377 31263
rect 29377 31229 29411 31263
rect 29411 31229 29420 31263
rect 29368 31220 29420 31229
rect 31760 31467 31812 31476
rect 31760 31433 31769 31467
rect 31769 31433 31803 31467
rect 31803 31433 31812 31467
rect 31760 31424 31812 31433
rect 32404 31424 32456 31476
rect 37556 31467 37608 31476
rect 37556 31433 37565 31467
rect 37565 31433 37599 31467
rect 37599 31433 37608 31467
rect 37556 31424 37608 31433
rect 38844 31424 38896 31476
rect 40408 31424 40460 31476
rect 47032 31467 47084 31476
rect 47032 31433 47041 31467
rect 47041 31433 47075 31467
rect 47075 31433 47084 31467
rect 47032 31424 47084 31433
rect 47124 31424 47176 31476
rect 32128 31356 32180 31408
rect 33968 31356 34020 31408
rect 32496 31331 32548 31340
rect 32496 31297 32505 31331
rect 32505 31297 32539 31331
rect 32539 31297 32548 31331
rect 32496 31288 32548 31297
rect 32128 31220 32180 31272
rect 35900 31288 35952 31340
rect 37464 31331 37516 31340
rect 37464 31297 37473 31331
rect 37473 31297 37507 31331
rect 37507 31297 37516 31331
rect 37464 31288 37516 31297
rect 39212 31356 39264 31408
rect 34060 31263 34112 31272
rect 34060 31229 34069 31263
rect 34069 31229 34103 31263
rect 34103 31229 34112 31263
rect 34060 31220 34112 31229
rect 33600 31152 33652 31204
rect 38660 31288 38712 31340
rect 38752 31331 38804 31340
rect 38752 31297 38761 31331
rect 38761 31297 38795 31331
rect 38795 31297 38804 31331
rect 38752 31288 38804 31297
rect 38936 31288 38988 31340
rect 40684 31288 40736 31340
rect 41604 31288 41656 31340
rect 46480 31288 46532 31340
rect 40592 31220 40644 31272
rect 41144 31263 41196 31272
rect 41144 31229 41153 31263
rect 41153 31229 41187 31263
rect 41187 31229 41196 31263
rect 41144 31220 41196 31229
rect 41328 31220 41380 31272
rect 42800 31220 42852 31272
rect 43536 31220 43588 31272
rect 38568 31152 38620 31204
rect 46940 31152 46992 31204
rect 27896 31127 27948 31136
rect 27896 31093 27905 31127
rect 27905 31093 27939 31127
rect 27939 31093 27948 31127
rect 27896 31084 27948 31093
rect 31208 31084 31260 31136
rect 32496 31084 32548 31136
rect 35440 31127 35492 31136
rect 35440 31093 35449 31127
rect 35449 31093 35483 31127
rect 35483 31093 35492 31127
rect 35440 31084 35492 31093
rect 35900 31127 35952 31136
rect 35900 31093 35909 31127
rect 35909 31093 35943 31127
rect 35943 31093 35952 31127
rect 35900 31084 35952 31093
rect 38108 31127 38160 31136
rect 38108 31093 38117 31127
rect 38117 31093 38151 31127
rect 38151 31093 38160 31127
rect 38108 31084 38160 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 30104 30923 30156 30932
rect 30104 30889 30113 30923
rect 30113 30889 30147 30923
rect 30147 30889 30156 30923
rect 30104 30880 30156 30889
rect 33600 30923 33652 30932
rect 33600 30889 33609 30923
rect 33609 30889 33643 30923
rect 33643 30889 33652 30923
rect 33600 30880 33652 30889
rect 40592 30880 40644 30932
rect 29736 30787 29788 30796
rect 29736 30753 29745 30787
rect 29745 30753 29779 30787
rect 29779 30753 29788 30787
rect 29736 30744 29788 30753
rect 31208 30787 31260 30796
rect 31208 30753 31217 30787
rect 31217 30753 31251 30787
rect 31251 30753 31260 30787
rect 31208 30744 31260 30753
rect 42340 30744 42392 30796
rect 44088 30880 44140 30932
rect 45836 30923 45888 30932
rect 45836 30889 45845 30923
rect 45845 30889 45879 30923
rect 45879 30889 45888 30923
rect 45836 30880 45888 30889
rect 43352 30812 43404 30864
rect 26516 30719 26568 30728
rect 26516 30685 26525 30719
rect 26525 30685 26559 30719
rect 26559 30685 26568 30719
rect 26516 30676 26568 30685
rect 26608 30719 26660 30728
rect 26608 30685 26617 30719
rect 26617 30685 26651 30719
rect 26651 30685 26660 30719
rect 26792 30719 26844 30728
rect 26608 30676 26660 30685
rect 26792 30685 26801 30719
rect 26801 30685 26835 30719
rect 26835 30685 26844 30719
rect 26792 30676 26844 30685
rect 27160 30676 27212 30728
rect 27436 30676 27488 30728
rect 30380 30676 30432 30728
rect 31392 30719 31444 30728
rect 31392 30685 31401 30719
rect 31401 30685 31435 30719
rect 31435 30685 31444 30719
rect 31392 30676 31444 30685
rect 32220 30719 32272 30728
rect 32220 30685 32229 30719
rect 32229 30685 32263 30719
rect 32263 30685 32272 30719
rect 32220 30676 32272 30685
rect 34060 30676 34112 30728
rect 37464 30719 37516 30728
rect 37464 30685 37473 30719
rect 37473 30685 37507 30719
rect 37507 30685 37516 30719
rect 37464 30676 37516 30685
rect 38108 30676 38160 30728
rect 40776 30719 40828 30728
rect 33140 30608 33192 30660
rect 35900 30608 35952 30660
rect 40776 30685 40785 30719
rect 40785 30685 40819 30719
rect 40819 30685 40828 30719
rect 40776 30676 40828 30685
rect 43536 30719 43588 30728
rect 41144 30608 41196 30660
rect 43536 30685 43545 30719
rect 43545 30685 43579 30719
rect 43579 30685 43588 30719
rect 43536 30676 43588 30685
rect 45560 30744 45612 30796
rect 45376 30719 45428 30728
rect 45376 30685 45383 30719
rect 45383 30685 45428 30719
rect 45376 30676 45428 30685
rect 45836 30676 45888 30728
rect 26608 30540 26660 30592
rect 31668 30540 31720 30592
rect 36176 30540 36228 30592
rect 40040 30540 40092 30592
rect 42892 30583 42944 30592
rect 42892 30549 42901 30583
rect 42901 30549 42935 30583
rect 42935 30549 42944 30583
rect 42892 30540 42944 30549
rect 43260 30540 43312 30592
rect 45192 30540 45244 30592
rect 46020 30540 46072 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 23480 30336 23532 30388
rect 26056 30336 26108 30388
rect 30012 30336 30064 30388
rect 33140 30379 33192 30388
rect 33140 30345 33149 30379
rect 33149 30345 33183 30379
rect 33183 30345 33192 30379
rect 33140 30336 33192 30345
rect 40776 30336 40828 30388
rect 41144 30379 41196 30388
rect 41144 30345 41153 30379
rect 41153 30345 41187 30379
rect 41187 30345 41196 30379
rect 41144 30336 41196 30345
rect 23296 30268 23348 30320
rect 31392 30268 31444 30320
rect 23388 30200 23440 30252
rect 31668 30243 31720 30252
rect 31668 30209 31677 30243
rect 31677 30209 31711 30243
rect 31711 30209 31720 30243
rect 31668 30200 31720 30209
rect 32128 30200 32180 30252
rect 32312 30243 32364 30252
rect 32312 30209 32321 30243
rect 32321 30209 32355 30243
rect 32355 30209 32364 30243
rect 32312 30200 32364 30209
rect 36176 30268 36228 30320
rect 35440 30200 35492 30252
rect 38844 30243 38896 30252
rect 38844 30209 38853 30243
rect 38853 30209 38887 30243
rect 38887 30209 38896 30243
rect 38844 30200 38896 30209
rect 40500 30268 40552 30320
rect 41328 30268 41380 30320
rect 39764 30243 39816 30252
rect 39764 30209 39773 30243
rect 39773 30209 39807 30243
rect 39807 30209 39816 30243
rect 39764 30200 39816 30209
rect 40224 30200 40276 30252
rect 40592 30243 40644 30252
rect 40592 30209 40601 30243
rect 40601 30209 40635 30243
rect 40635 30209 40644 30243
rect 40592 30200 40644 30209
rect 40776 30243 40828 30252
rect 40776 30209 40785 30243
rect 40785 30209 40819 30243
rect 40819 30209 40828 30243
rect 40776 30200 40828 30209
rect 41972 30200 42024 30252
rect 42892 30268 42944 30320
rect 43076 30200 43128 30252
rect 45008 30243 45060 30252
rect 45008 30209 45017 30243
rect 45017 30209 45051 30243
rect 45051 30209 45060 30243
rect 45008 30200 45060 30209
rect 45376 30243 45428 30252
rect 45376 30209 45385 30243
rect 45385 30209 45419 30243
rect 45419 30209 45428 30243
rect 45376 30200 45428 30209
rect 42892 30132 42944 30184
rect 45100 30175 45152 30184
rect 45100 30141 45109 30175
rect 45109 30141 45143 30175
rect 45143 30141 45152 30175
rect 45100 30132 45152 30141
rect 45192 30175 45244 30184
rect 45192 30141 45201 30175
rect 45201 30141 45235 30175
rect 45235 30141 45244 30175
rect 45836 30200 45888 30252
rect 47492 30200 47544 30252
rect 47676 30200 47728 30252
rect 45192 30132 45244 30141
rect 46204 30132 46256 30184
rect 44088 30064 44140 30116
rect 24400 29996 24452 30048
rect 31576 29996 31628 30048
rect 35348 30039 35400 30048
rect 35348 30005 35357 30039
rect 35357 30005 35391 30039
rect 35391 30005 35400 30039
rect 35348 29996 35400 30005
rect 38936 30039 38988 30048
rect 38936 30005 38945 30039
rect 38945 30005 38979 30039
rect 38979 30005 38988 30039
rect 38936 29996 38988 30005
rect 43628 29996 43680 30048
rect 45560 30039 45612 30048
rect 45560 30005 45569 30039
rect 45569 30005 45603 30039
rect 45603 30005 45612 30039
rect 45560 29996 45612 30005
rect 46020 29996 46072 30048
rect 47216 30039 47268 30048
rect 47216 30005 47225 30039
rect 47225 30005 47259 30039
rect 47259 30005 47268 30039
rect 47216 29996 47268 30005
rect 47860 30039 47912 30048
rect 47860 30005 47869 30039
rect 47869 30005 47903 30039
rect 47903 30005 47912 30039
rect 47860 29996 47912 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 23388 29835 23440 29844
rect 23388 29801 23397 29835
rect 23397 29801 23431 29835
rect 23431 29801 23440 29835
rect 23388 29792 23440 29801
rect 27436 29792 27488 29844
rect 32312 29792 32364 29844
rect 39764 29792 39816 29844
rect 40040 29835 40092 29844
rect 40040 29801 40049 29835
rect 40049 29801 40083 29835
rect 40083 29801 40092 29835
rect 40040 29792 40092 29801
rect 40776 29792 40828 29844
rect 45192 29792 45244 29844
rect 24768 29724 24820 29776
rect 23296 29588 23348 29640
rect 23572 29588 23624 29640
rect 24400 29656 24452 29708
rect 35440 29724 35492 29776
rect 24032 29631 24084 29640
rect 24032 29597 24041 29631
rect 24041 29597 24075 29631
rect 24075 29597 24084 29631
rect 24032 29588 24084 29597
rect 26608 29631 26660 29640
rect 26608 29597 26617 29631
rect 26617 29597 26651 29631
rect 26651 29597 26660 29631
rect 26608 29588 26660 29597
rect 28724 29588 28776 29640
rect 31576 29631 31628 29640
rect 31576 29597 31610 29631
rect 31610 29597 31628 29631
rect 26424 29520 26476 29572
rect 23940 29452 23992 29504
rect 24584 29452 24636 29504
rect 26516 29495 26568 29504
rect 26516 29461 26525 29495
rect 26525 29461 26559 29495
rect 26559 29461 26568 29495
rect 26516 29452 26568 29461
rect 27160 29520 27212 29572
rect 27896 29452 27948 29504
rect 31576 29588 31628 29597
rect 34244 29588 34296 29640
rect 38844 29656 38896 29708
rect 36176 29631 36228 29640
rect 36176 29597 36185 29631
rect 36185 29597 36219 29631
rect 36219 29597 36228 29631
rect 36176 29588 36228 29597
rect 38936 29631 38988 29640
rect 38936 29597 38945 29631
rect 38945 29597 38979 29631
rect 38979 29597 38988 29631
rect 38936 29588 38988 29597
rect 41328 29656 41380 29708
rect 40224 29631 40276 29640
rect 40224 29597 40233 29631
rect 40233 29597 40267 29631
rect 40267 29597 40276 29631
rect 40224 29588 40276 29597
rect 40500 29588 40552 29640
rect 40592 29631 40644 29640
rect 40592 29597 40601 29631
rect 40601 29597 40635 29631
rect 40635 29597 40644 29631
rect 40592 29588 40644 29597
rect 41972 29588 42024 29640
rect 47216 29656 47268 29708
rect 43628 29588 43680 29640
rect 43720 29631 43772 29640
rect 43720 29597 43729 29631
rect 43729 29597 43763 29631
rect 43763 29597 43772 29631
rect 43720 29588 43772 29597
rect 43996 29588 44048 29640
rect 45008 29588 45060 29640
rect 45744 29588 45796 29640
rect 34612 29520 34664 29572
rect 35624 29520 35676 29572
rect 45100 29520 45152 29572
rect 47860 29520 47912 29572
rect 48320 29563 48372 29572
rect 48320 29529 48329 29563
rect 48329 29529 48363 29563
rect 48363 29529 48372 29563
rect 48320 29520 48372 29529
rect 31760 29452 31812 29504
rect 32220 29452 32272 29504
rect 35900 29452 35952 29504
rect 36360 29495 36412 29504
rect 36360 29461 36369 29495
rect 36369 29461 36403 29495
rect 36403 29461 36412 29495
rect 36360 29452 36412 29461
rect 43260 29452 43312 29504
rect 44088 29495 44140 29504
rect 44088 29461 44097 29495
rect 44097 29461 44131 29495
rect 44131 29461 44140 29495
rect 44088 29452 44140 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 23296 29291 23348 29300
rect 23296 29257 23305 29291
rect 23305 29257 23339 29291
rect 23339 29257 23348 29291
rect 23296 29248 23348 29257
rect 23940 29291 23992 29300
rect 23940 29257 23949 29291
rect 23949 29257 23983 29291
rect 23983 29257 23992 29291
rect 23940 29248 23992 29257
rect 24032 29248 24084 29300
rect 27160 29291 27212 29300
rect 24676 29180 24728 29232
rect 27160 29257 27169 29291
rect 27169 29257 27203 29291
rect 27203 29257 27212 29291
rect 27160 29248 27212 29257
rect 24584 29155 24636 29164
rect 24584 29121 24593 29155
rect 24593 29121 24627 29155
rect 24627 29121 24636 29155
rect 24584 29112 24636 29121
rect 26424 29155 26476 29164
rect 26424 29121 26433 29155
rect 26433 29121 26467 29155
rect 26467 29121 26476 29155
rect 26424 29112 26476 29121
rect 26608 29155 26660 29164
rect 26608 29121 26617 29155
rect 26617 29121 26651 29155
rect 26651 29121 26660 29155
rect 26608 29112 26660 29121
rect 27436 29155 27488 29164
rect 27436 29121 27445 29155
rect 27445 29121 27479 29155
rect 27479 29121 27488 29155
rect 27436 29112 27488 29121
rect 23664 29087 23716 29096
rect 23664 29053 23673 29087
rect 23673 29053 23707 29087
rect 23707 29053 23716 29087
rect 23664 29044 23716 29053
rect 24768 29044 24820 29096
rect 27620 29155 27672 29164
rect 27620 29121 27629 29155
rect 27629 29121 27663 29155
rect 27663 29121 27672 29155
rect 29368 29180 29420 29232
rect 29828 29180 29880 29232
rect 33416 29180 33468 29232
rect 34244 29223 34296 29232
rect 34244 29189 34253 29223
rect 34253 29189 34287 29223
rect 34287 29189 34296 29223
rect 35716 29248 35768 29300
rect 40224 29248 40276 29300
rect 40776 29291 40828 29300
rect 40776 29257 40785 29291
rect 40785 29257 40819 29291
rect 40819 29257 40828 29291
rect 40776 29248 40828 29257
rect 41972 29291 42024 29300
rect 41972 29257 41981 29291
rect 41981 29257 42015 29291
rect 42015 29257 42024 29291
rect 41972 29248 42024 29257
rect 43076 29248 43128 29300
rect 43260 29291 43312 29300
rect 43260 29257 43269 29291
rect 43269 29257 43303 29291
rect 43303 29257 43312 29291
rect 43260 29248 43312 29257
rect 43720 29248 43772 29300
rect 34244 29180 34296 29189
rect 27620 29112 27672 29121
rect 28724 29155 28776 29164
rect 28724 29121 28733 29155
rect 28733 29121 28767 29155
rect 28767 29121 28776 29155
rect 28724 29112 28776 29121
rect 30748 29155 30800 29164
rect 30748 29121 30757 29155
rect 30757 29121 30791 29155
rect 30791 29121 30800 29155
rect 30748 29112 30800 29121
rect 35348 29155 35400 29164
rect 35348 29121 35357 29155
rect 35357 29121 35391 29155
rect 35391 29121 35400 29155
rect 35348 29112 35400 29121
rect 24492 28951 24544 28960
rect 24492 28917 24501 28951
rect 24501 28917 24535 28951
rect 24535 28917 24544 28951
rect 24492 28908 24544 28917
rect 26792 28908 26844 28960
rect 29920 29044 29972 29096
rect 27896 28908 27948 28960
rect 34612 29019 34664 29028
rect 34612 28985 34621 29019
rect 34621 28985 34655 29019
rect 34655 28985 34664 29019
rect 34612 28976 34664 28985
rect 29920 28908 29972 28960
rect 34704 28951 34756 28960
rect 34704 28917 34713 28951
rect 34713 28917 34747 28951
rect 34747 28917 34756 28951
rect 34704 28908 34756 28917
rect 35256 28908 35308 28960
rect 35992 29112 36044 29164
rect 38752 29180 38804 29232
rect 38016 29112 38068 29164
rect 40684 29155 40736 29164
rect 35900 29044 35952 29096
rect 37464 29087 37516 29096
rect 37464 29053 37473 29087
rect 37473 29053 37507 29087
rect 37507 29053 37516 29087
rect 37464 29044 37516 29053
rect 40684 29121 40693 29155
rect 40693 29121 40727 29155
rect 40727 29121 40736 29155
rect 40684 29112 40736 29121
rect 41512 29112 41564 29164
rect 44088 29180 44140 29232
rect 40224 29044 40276 29096
rect 42340 29044 42392 29096
rect 43904 29112 43956 29164
rect 45652 29112 45704 29164
rect 45560 29087 45612 29096
rect 45560 29053 45569 29087
rect 45569 29053 45603 29087
rect 45603 29053 45612 29087
rect 45560 29044 45612 29053
rect 36636 28951 36688 28960
rect 36636 28917 36645 28951
rect 36645 28917 36679 28951
rect 36679 28917 36688 28951
rect 36636 28908 36688 28917
rect 38936 28976 38988 29028
rect 40408 28976 40460 29028
rect 38476 28908 38528 28960
rect 45836 28908 45888 28960
rect 47952 28951 48004 28960
rect 47952 28917 47961 28951
rect 47961 28917 47995 28951
rect 47995 28917 48004 28951
rect 47952 28908 48004 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 23664 28704 23716 28756
rect 26608 28704 26660 28756
rect 27620 28704 27672 28756
rect 30748 28704 30800 28756
rect 26700 28636 26752 28688
rect 23664 28568 23716 28620
rect 24584 28568 24636 28620
rect 26792 28611 26844 28620
rect 24492 28500 24544 28552
rect 26792 28577 26801 28611
rect 26801 28577 26835 28611
rect 26835 28577 26844 28611
rect 26792 28568 26844 28577
rect 22652 28364 22704 28416
rect 23388 28407 23440 28416
rect 23388 28373 23397 28407
rect 23397 28373 23431 28407
rect 23431 28373 23440 28407
rect 23388 28364 23440 28373
rect 24676 28432 24728 28484
rect 24952 28364 25004 28416
rect 26516 28500 26568 28552
rect 27896 28543 27948 28552
rect 27896 28509 27905 28543
rect 27905 28509 27939 28543
rect 27939 28509 27948 28543
rect 27896 28500 27948 28509
rect 30012 28543 30064 28552
rect 30012 28509 30021 28543
rect 30021 28509 30055 28543
rect 30055 28509 30064 28543
rect 30012 28500 30064 28509
rect 31760 28500 31812 28552
rect 35992 28704 36044 28756
rect 36912 28704 36964 28756
rect 43996 28704 44048 28756
rect 45652 28704 45704 28756
rect 35440 28611 35492 28620
rect 27436 28432 27488 28484
rect 30656 28432 30708 28484
rect 32956 28432 33008 28484
rect 34704 28432 34756 28484
rect 35440 28577 35449 28611
rect 35449 28577 35483 28611
rect 35483 28577 35492 28611
rect 35440 28568 35492 28577
rect 36360 28636 36412 28688
rect 39212 28636 39264 28688
rect 35624 28500 35676 28552
rect 35992 28568 36044 28620
rect 35900 28500 35952 28552
rect 36636 28500 36688 28552
rect 40132 28568 40184 28620
rect 40684 28568 40736 28620
rect 41144 28568 41196 28620
rect 46848 28636 46900 28688
rect 45836 28568 45888 28620
rect 47952 28568 48004 28620
rect 48228 28611 48280 28620
rect 48228 28577 48237 28611
rect 48237 28577 48271 28611
rect 48271 28577 48280 28611
rect 48228 28568 48280 28577
rect 40224 28543 40276 28552
rect 40224 28509 40233 28543
rect 40233 28509 40267 28543
rect 40267 28509 40276 28543
rect 40224 28500 40276 28509
rect 40408 28500 40460 28552
rect 41512 28543 41564 28552
rect 41512 28509 41521 28543
rect 41521 28509 41555 28543
rect 41555 28509 41564 28543
rect 41512 28500 41564 28509
rect 41604 28543 41656 28552
rect 41604 28509 41613 28543
rect 41613 28509 41647 28543
rect 41647 28509 41656 28543
rect 41604 28500 41656 28509
rect 42432 28543 42484 28552
rect 42432 28509 42441 28543
rect 42441 28509 42475 28543
rect 42475 28509 42484 28543
rect 42432 28500 42484 28509
rect 43812 28500 43864 28552
rect 45744 28543 45796 28552
rect 45744 28509 45753 28543
rect 45753 28509 45787 28543
rect 45787 28509 45796 28543
rect 45744 28500 45796 28509
rect 45928 28543 45980 28552
rect 45928 28509 45937 28543
rect 45937 28509 45971 28543
rect 45971 28509 45980 28543
rect 45928 28500 45980 28509
rect 47860 28432 47912 28484
rect 26608 28364 26660 28416
rect 29920 28407 29972 28416
rect 29920 28373 29929 28407
rect 29929 28373 29963 28407
rect 29963 28373 29972 28407
rect 29920 28364 29972 28373
rect 32312 28364 32364 28416
rect 35532 28364 35584 28416
rect 36268 28364 36320 28416
rect 42340 28407 42392 28416
rect 42340 28373 42349 28407
rect 42349 28373 42383 28407
rect 42383 28373 42392 28407
rect 42340 28364 42392 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 12992 28160 13044 28212
rect 23388 28092 23440 28144
rect 24952 28092 25004 28144
rect 25596 28092 25648 28144
rect 26332 28092 26384 28144
rect 26608 28135 26660 28144
rect 26608 28101 26617 28135
rect 26617 28101 26651 28135
rect 26651 28101 26660 28135
rect 26608 28092 26660 28101
rect 32956 28160 33008 28212
rect 38016 28203 38068 28212
rect 38016 28169 38025 28203
rect 38025 28169 38059 28203
rect 38059 28169 38068 28203
rect 38016 28160 38068 28169
rect 22928 28067 22980 28076
rect 22928 28033 22937 28067
rect 22937 28033 22971 28067
rect 22971 28033 22980 28067
rect 22928 28024 22980 28033
rect 23204 28067 23256 28076
rect 23204 28033 23213 28067
rect 23213 28033 23247 28067
rect 23247 28033 23256 28067
rect 23204 28024 23256 28033
rect 23664 28067 23716 28076
rect 23664 28033 23673 28067
rect 23673 28033 23707 28067
rect 23707 28033 23716 28067
rect 23664 28024 23716 28033
rect 23848 28067 23900 28076
rect 23848 28033 23857 28067
rect 23857 28033 23891 28067
rect 23891 28033 23900 28067
rect 23848 28024 23900 28033
rect 24124 28024 24176 28076
rect 23020 27956 23072 28008
rect 23756 27888 23808 27940
rect 26516 28024 26568 28076
rect 29920 28024 29972 28076
rect 30656 28024 30708 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 24492 27956 24544 28008
rect 24768 27888 24820 27940
rect 25228 27931 25280 27940
rect 25228 27897 25237 27931
rect 25237 27897 25271 27931
rect 25271 27897 25280 27931
rect 25228 27888 25280 27897
rect 23480 27820 23532 27872
rect 24860 27820 24912 27872
rect 32588 27999 32640 28008
rect 32588 27965 32597 27999
rect 32597 27965 32631 27999
rect 32631 27965 32640 27999
rect 32588 27956 32640 27965
rect 32680 27956 32732 28008
rect 28540 27820 28592 27872
rect 30380 27820 30432 27872
rect 31944 27820 31996 27872
rect 34796 27820 34848 27872
rect 36360 28092 36412 28144
rect 38936 28160 38988 28212
rect 40132 28160 40184 28212
rect 41512 28160 41564 28212
rect 45744 28203 45796 28212
rect 45744 28169 45759 28203
rect 45759 28169 45793 28203
rect 45793 28169 45796 28203
rect 47860 28203 47912 28212
rect 45744 28160 45796 28169
rect 47860 28169 47869 28203
rect 47869 28169 47903 28203
rect 47903 28169 47912 28203
rect 47860 28160 47912 28169
rect 35992 28024 36044 28076
rect 38476 28092 38528 28144
rect 38016 28024 38068 28076
rect 39120 28024 39172 28076
rect 42340 28092 42392 28144
rect 45836 28135 45888 28144
rect 35440 27956 35492 28008
rect 38476 27956 38528 28008
rect 35624 27888 35676 27940
rect 43168 28067 43220 28076
rect 43168 28033 43202 28067
rect 43202 28033 43220 28067
rect 43168 28024 43220 28033
rect 42892 27999 42944 28008
rect 42892 27965 42901 27999
rect 42901 27965 42935 27999
rect 42935 27965 42944 27999
rect 42892 27956 42944 27965
rect 45836 28101 45845 28135
rect 45845 28101 45879 28135
rect 45879 28101 45888 28135
rect 45836 28092 45888 28101
rect 45744 28024 45796 28076
rect 45928 28067 45980 28076
rect 45928 28033 45937 28067
rect 45937 28033 45971 28067
rect 45971 28033 45980 28067
rect 45928 28024 45980 28033
rect 46480 28024 46532 28076
rect 47492 28024 47544 28076
rect 43812 27820 43864 27872
rect 46388 27863 46440 27872
rect 46388 27829 46397 27863
rect 46397 27829 46431 27863
rect 46431 27829 46440 27863
rect 46388 27820 46440 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 22928 27616 22980 27668
rect 26608 27616 26660 27668
rect 39120 27659 39172 27668
rect 39120 27625 39129 27659
rect 39129 27625 39163 27659
rect 39163 27625 39172 27659
rect 39120 27616 39172 27625
rect 40224 27659 40276 27668
rect 40224 27625 40233 27659
rect 40233 27625 40267 27659
rect 40267 27625 40276 27659
rect 40224 27616 40276 27625
rect 23020 27548 23072 27600
rect 24584 27548 24636 27600
rect 25596 27548 25648 27600
rect 32680 27548 32732 27600
rect 33784 27548 33836 27600
rect 38016 27548 38068 27600
rect 39212 27591 39264 27600
rect 39212 27557 39221 27591
rect 39221 27557 39255 27591
rect 39255 27557 39264 27591
rect 39212 27548 39264 27557
rect 23572 27523 23624 27532
rect 23572 27489 23581 27523
rect 23581 27489 23615 27523
rect 23615 27489 23624 27523
rect 23572 27480 23624 27489
rect 23756 27523 23808 27532
rect 23756 27489 23765 27523
rect 23765 27489 23799 27523
rect 23799 27489 23808 27523
rect 23756 27480 23808 27489
rect 22652 27455 22704 27464
rect 22652 27421 22661 27455
rect 22661 27421 22695 27455
rect 22695 27421 22704 27455
rect 22652 27412 22704 27421
rect 23112 27412 23164 27464
rect 26332 27480 26384 27532
rect 29828 27480 29880 27532
rect 31852 27480 31904 27532
rect 32312 27480 32364 27532
rect 24400 27412 24452 27464
rect 24860 27455 24912 27464
rect 24860 27421 24894 27455
rect 24894 27421 24912 27455
rect 24860 27412 24912 27421
rect 26608 27455 26660 27464
rect 26608 27421 26617 27455
rect 26617 27421 26651 27455
rect 26651 27421 26660 27455
rect 26608 27412 26660 27421
rect 25596 27344 25648 27396
rect 25688 27344 25740 27396
rect 27528 27412 27580 27464
rect 31944 27455 31996 27464
rect 31944 27421 31953 27455
rect 31953 27421 31987 27455
rect 31987 27421 31996 27455
rect 31944 27412 31996 27421
rect 35532 27480 35584 27532
rect 40316 27548 40368 27600
rect 41604 27616 41656 27668
rect 42432 27616 42484 27668
rect 43168 27659 43220 27668
rect 43168 27625 43177 27659
rect 43177 27625 43211 27659
rect 43211 27625 43220 27659
rect 43168 27616 43220 27625
rect 43904 27659 43956 27668
rect 43904 27625 43913 27659
rect 43913 27625 43947 27659
rect 43947 27625 43956 27659
rect 43904 27616 43956 27625
rect 45928 27616 45980 27668
rect 46480 27616 46532 27668
rect 42892 27548 42944 27600
rect 43260 27548 43312 27600
rect 45560 27548 45612 27600
rect 35348 27455 35400 27464
rect 35348 27421 35357 27455
rect 35357 27421 35391 27455
rect 35391 27421 35400 27455
rect 35348 27412 35400 27421
rect 41512 27480 41564 27532
rect 40316 27412 40368 27464
rect 41604 27412 41656 27464
rect 43352 27412 43404 27464
rect 30196 27387 30248 27396
rect 30196 27353 30230 27387
rect 30230 27353 30248 27387
rect 33692 27387 33744 27396
rect 30196 27344 30248 27353
rect 33692 27353 33701 27387
rect 33701 27353 33735 27387
rect 33735 27353 33744 27387
rect 33692 27344 33744 27353
rect 35900 27344 35952 27396
rect 40132 27344 40184 27396
rect 41052 27344 41104 27396
rect 43720 27387 43772 27396
rect 43720 27353 43729 27387
rect 43729 27353 43763 27387
rect 43763 27353 43772 27387
rect 43720 27344 43772 27353
rect 23296 27319 23348 27328
rect 23296 27285 23305 27319
rect 23305 27285 23339 27319
rect 23339 27285 23348 27319
rect 23296 27276 23348 27285
rect 25964 27319 26016 27328
rect 25964 27285 25973 27319
rect 25973 27285 26007 27319
rect 26007 27285 26016 27319
rect 25964 27276 26016 27285
rect 27620 27276 27672 27328
rect 28172 27319 28224 27328
rect 28172 27285 28181 27319
rect 28181 27285 28215 27319
rect 28215 27285 28224 27319
rect 28172 27276 28224 27285
rect 30656 27276 30708 27328
rect 33784 27319 33836 27328
rect 33784 27285 33793 27319
rect 33793 27285 33827 27319
rect 33827 27285 33836 27319
rect 33784 27276 33836 27285
rect 35348 27276 35400 27328
rect 40408 27276 40460 27328
rect 42432 27276 42484 27328
rect 43628 27276 43680 27328
rect 45652 27480 45704 27532
rect 46848 27523 46900 27532
rect 46848 27489 46857 27523
rect 46857 27489 46891 27523
rect 46891 27489 46900 27523
rect 46848 27480 46900 27489
rect 46756 27412 46808 27464
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 23388 27115 23440 27124
rect 23388 27081 23397 27115
rect 23397 27081 23431 27115
rect 23431 27081 23440 27115
rect 23388 27072 23440 27081
rect 26608 27072 26660 27124
rect 22928 26936 22980 26988
rect 23480 26979 23532 26988
rect 23480 26945 23489 26979
rect 23489 26945 23523 26979
rect 23523 26945 23532 26979
rect 25688 27004 25740 27056
rect 30196 27072 30248 27124
rect 31024 27115 31076 27124
rect 23480 26936 23532 26945
rect 23204 26868 23256 26920
rect 24768 26868 24820 26920
rect 25964 26936 26016 26988
rect 27436 26979 27488 26988
rect 26332 26868 26384 26920
rect 27436 26945 27445 26979
rect 27445 26945 27479 26979
rect 27479 26945 27488 26979
rect 27436 26936 27488 26945
rect 27528 26979 27580 26988
rect 27528 26945 27538 26979
rect 27538 26945 27572 26979
rect 27572 26945 27580 26979
rect 27804 26979 27856 26988
rect 27528 26936 27580 26945
rect 27804 26945 27813 26979
rect 27813 26945 27847 26979
rect 27847 26945 27856 26979
rect 27804 26936 27856 26945
rect 30380 27004 30432 27056
rect 31024 27081 31033 27115
rect 31033 27081 31067 27115
rect 31067 27081 31076 27115
rect 31024 27072 31076 27081
rect 30656 27047 30708 27056
rect 30656 27013 30665 27047
rect 30665 27013 30699 27047
rect 30699 27013 30708 27047
rect 30656 27004 30708 27013
rect 31300 27004 31352 27056
rect 31944 27072 31996 27124
rect 35348 27072 35400 27124
rect 36912 27115 36964 27124
rect 36912 27081 36921 27115
rect 36921 27081 36955 27115
rect 36955 27081 36964 27115
rect 36912 27072 36964 27081
rect 43904 27072 43956 27124
rect 46756 27072 46808 27124
rect 33508 26936 33560 26988
rect 33692 26936 33744 26988
rect 35072 26979 35124 26988
rect 32956 26911 33008 26920
rect 32956 26877 32965 26911
rect 32965 26877 32999 26911
rect 32999 26877 33008 26911
rect 32956 26868 33008 26877
rect 35072 26945 35081 26979
rect 35081 26945 35115 26979
rect 35115 26945 35124 26979
rect 35072 26936 35124 26945
rect 38292 27004 38344 27056
rect 43720 27004 43772 27056
rect 46388 27004 46440 27056
rect 36176 26936 36228 26988
rect 43628 26979 43680 26988
rect 43628 26945 43637 26979
rect 43637 26945 43671 26979
rect 43671 26945 43680 26979
rect 43628 26936 43680 26945
rect 45560 26936 45612 26988
rect 46940 26936 46992 26988
rect 47584 26936 47636 26988
rect 27344 26800 27396 26852
rect 30656 26800 30708 26852
rect 23572 26732 23624 26784
rect 24676 26732 24728 26784
rect 27436 26732 27488 26784
rect 27712 26775 27764 26784
rect 27712 26741 27721 26775
rect 27721 26741 27755 26775
rect 27755 26741 27764 26775
rect 31852 26800 31904 26852
rect 36728 26800 36780 26852
rect 37188 26800 37240 26852
rect 41604 26800 41656 26852
rect 43352 26843 43404 26852
rect 43352 26809 43361 26843
rect 43361 26809 43395 26843
rect 43395 26809 43404 26843
rect 43352 26800 43404 26809
rect 27712 26732 27764 26741
rect 34796 26775 34848 26784
rect 34796 26741 34805 26775
rect 34805 26741 34839 26775
rect 34839 26741 34848 26775
rect 34796 26732 34848 26741
rect 35072 26732 35124 26784
rect 37832 26732 37884 26784
rect 38292 26732 38344 26784
rect 45652 26732 45704 26784
rect 47860 26775 47912 26784
rect 47860 26741 47869 26775
rect 47869 26741 47903 26775
rect 47903 26741 47912 26775
rect 47860 26732 47912 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 31760 26528 31812 26580
rect 32956 26528 33008 26580
rect 33508 26571 33560 26580
rect 33508 26537 33517 26571
rect 33517 26537 33551 26571
rect 33551 26537 33560 26571
rect 33508 26528 33560 26537
rect 36544 26528 36596 26580
rect 39488 26528 39540 26580
rect 40408 26571 40460 26580
rect 40408 26537 40417 26571
rect 40417 26537 40451 26571
rect 40451 26537 40460 26571
rect 40408 26528 40460 26537
rect 43628 26528 43680 26580
rect 37188 26460 37240 26512
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 26332 26324 26384 26333
rect 28080 26392 28132 26444
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 27712 26324 27764 26376
rect 27804 26324 27856 26376
rect 34796 26392 34848 26444
rect 35440 26435 35492 26444
rect 35440 26401 35449 26435
rect 35449 26401 35483 26435
rect 35483 26401 35492 26435
rect 35440 26392 35492 26401
rect 40224 26460 40276 26512
rect 35348 26367 35400 26376
rect 35348 26333 35357 26367
rect 35357 26333 35391 26367
rect 35391 26333 35400 26367
rect 35348 26324 35400 26333
rect 38016 26367 38068 26376
rect 38016 26333 38025 26367
rect 38025 26333 38059 26367
rect 38059 26333 38068 26367
rect 38016 26324 38068 26333
rect 38476 26324 38528 26376
rect 39488 26367 39540 26376
rect 39488 26333 39497 26367
rect 39497 26333 39531 26367
rect 39531 26333 39540 26367
rect 39488 26324 39540 26333
rect 43904 26367 43956 26376
rect 43904 26333 43913 26367
rect 43913 26333 43947 26367
rect 43947 26333 43956 26367
rect 44548 26367 44600 26376
rect 43904 26324 43956 26333
rect 44548 26333 44557 26367
rect 44557 26333 44591 26367
rect 44591 26333 44600 26367
rect 44548 26324 44600 26333
rect 47860 26392 47912 26444
rect 48228 26435 48280 26444
rect 48228 26401 48237 26435
rect 48237 26401 48271 26435
rect 48271 26401 48280 26435
rect 48228 26392 48280 26401
rect 31208 26299 31260 26308
rect 31208 26265 31217 26299
rect 31217 26265 31251 26299
rect 31251 26265 31260 26299
rect 31208 26256 31260 26265
rect 36728 26256 36780 26308
rect 36820 26256 36872 26308
rect 38752 26256 38804 26308
rect 45652 26256 45704 26308
rect 47952 26256 48004 26308
rect 27344 26188 27396 26240
rect 27804 26231 27856 26240
rect 27804 26197 27813 26231
rect 27813 26197 27847 26231
rect 27847 26197 27856 26231
rect 27804 26188 27856 26197
rect 32588 26188 32640 26240
rect 37924 26188 37976 26240
rect 38660 26188 38712 26240
rect 40132 26188 40184 26240
rect 40224 26188 40276 26240
rect 43536 26188 43588 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 29828 25984 29880 26036
rect 35440 25984 35492 26036
rect 36176 26027 36228 26036
rect 36176 25993 36185 26027
rect 36185 25993 36219 26027
rect 36219 25993 36228 26027
rect 36176 25984 36228 25993
rect 36544 25984 36596 26036
rect 23388 25848 23440 25900
rect 27804 25916 27856 25968
rect 31208 25916 31260 25968
rect 27344 25891 27396 25900
rect 27344 25857 27353 25891
rect 27353 25857 27387 25891
rect 27387 25857 27396 25891
rect 27344 25848 27396 25857
rect 27988 25848 28040 25900
rect 30932 25848 30984 25900
rect 33692 25916 33744 25968
rect 35532 25891 35584 25900
rect 23940 25780 23992 25832
rect 22928 25712 22980 25764
rect 1584 25644 1636 25696
rect 22376 25644 22428 25696
rect 26332 25780 26384 25832
rect 24400 25644 24452 25696
rect 25412 25687 25464 25696
rect 25412 25653 25421 25687
rect 25421 25653 25455 25687
rect 25455 25653 25464 25687
rect 25412 25644 25464 25653
rect 27436 25644 27488 25696
rect 30748 25780 30800 25832
rect 35532 25857 35541 25891
rect 35541 25857 35575 25891
rect 35575 25857 35584 25891
rect 35532 25848 35584 25857
rect 36360 25848 36412 25900
rect 36728 25848 36780 25900
rect 37188 25848 37240 25900
rect 40224 25984 40276 26036
rect 44548 25984 44600 26036
rect 47216 25959 47268 25968
rect 36912 25780 36964 25832
rect 37832 25848 37884 25900
rect 40132 25848 40184 25900
rect 47216 25925 47225 25959
rect 47225 25925 47259 25959
rect 47259 25925 47268 25959
rect 47216 25916 47268 25925
rect 43260 25891 43312 25900
rect 43260 25857 43269 25891
rect 43269 25857 43303 25891
rect 43303 25857 43312 25891
rect 43260 25848 43312 25857
rect 43536 25891 43588 25900
rect 43536 25857 43570 25891
rect 43570 25857 43588 25891
rect 43536 25848 43588 25857
rect 47952 25891 48004 25900
rect 47952 25857 47961 25891
rect 47961 25857 47995 25891
rect 47995 25857 48004 25891
rect 47952 25848 48004 25857
rect 47124 25780 47176 25832
rect 46848 25712 46900 25764
rect 27712 25644 27764 25696
rect 30840 25687 30892 25696
rect 30840 25653 30849 25687
rect 30849 25653 30883 25687
rect 30883 25653 30892 25687
rect 30840 25644 30892 25653
rect 32496 25687 32548 25696
rect 32496 25653 32505 25687
rect 32505 25653 32539 25687
rect 32539 25653 32548 25687
rect 32496 25644 32548 25653
rect 38200 25644 38252 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 23388 25483 23440 25492
rect 23388 25449 23397 25483
rect 23397 25449 23431 25483
rect 23431 25449 23440 25483
rect 23388 25440 23440 25449
rect 23940 25440 23992 25492
rect 26332 25440 26384 25492
rect 28080 25483 28132 25492
rect 28080 25449 28089 25483
rect 28089 25449 28123 25483
rect 28123 25449 28132 25483
rect 28080 25440 28132 25449
rect 36360 25483 36412 25492
rect 36360 25449 36369 25483
rect 36369 25449 36403 25483
rect 36403 25449 36412 25483
rect 36360 25440 36412 25449
rect 38844 25372 38896 25424
rect 42248 25372 42300 25424
rect 46020 25372 46072 25424
rect 1584 25347 1636 25356
rect 1584 25313 1593 25347
rect 1593 25313 1627 25347
rect 1627 25313 1636 25347
rect 1584 25304 1636 25313
rect 2780 25347 2832 25356
rect 2780 25313 2789 25347
rect 2789 25313 2823 25347
rect 2823 25313 2832 25347
rect 2780 25304 2832 25313
rect 22744 25279 22796 25288
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 23296 25236 23348 25288
rect 1768 25211 1820 25220
rect 1768 25177 1777 25211
rect 1777 25177 1811 25211
rect 1811 25177 1820 25211
rect 1768 25168 1820 25177
rect 22376 25168 22428 25220
rect 23848 25279 23900 25288
rect 23848 25245 23857 25279
rect 23857 25245 23891 25279
rect 23891 25245 23900 25279
rect 23848 25236 23900 25245
rect 24032 25279 24084 25288
rect 24032 25245 24041 25279
rect 24041 25245 24075 25279
rect 24075 25245 24084 25279
rect 24032 25236 24084 25245
rect 24952 25236 25004 25288
rect 25412 25236 25464 25288
rect 28172 25304 28224 25356
rect 30932 25304 30984 25356
rect 32588 25304 32640 25356
rect 35348 25304 35400 25356
rect 24124 25168 24176 25220
rect 25320 25168 25372 25220
rect 22928 25143 22980 25152
rect 22928 25109 22937 25143
rect 22937 25109 22971 25143
rect 22971 25109 22980 25143
rect 22928 25100 22980 25109
rect 27896 25279 27948 25288
rect 27896 25245 27910 25279
rect 27910 25245 27944 25279
rect 27944 25245 27948 25279
rect 27896 25236 27948 25245
rect 31576 25279 31628 25288
rect 27620 25100 27672 25152
rect 27804 25211 27856 25220
rect 27804 25177 27813 25211
rect 27813 25177 27847 25211
rect 27847 25177 27856 25211
rect 27804 25168 27856 25177
rect 29828 25168 29880 25220
rect 31576 25245 31585 25279
rect 31585 25245 31619 25279
rect 31619 25245 31628 25279
rect 31576 25236 31628 25245
rect 36176 25236 36228 25288
rect 36912 25236 36964 25288
rect 39028 25279 39080 25288
rect 31760 25168 31812 25220
rect 35624 25168 35676 25220
rect 36268 25168 36320 25220
rect 39028 25245 39037 25279
rect 39037 25245 39071 25279
rect 39071 25245 39080 25279
rect 39028 25236 39080 25245
rect 42156 25279 42208 25288
rect 38752 25211 38804 25220
rect 38752 25177 38761 25211
rect 38761 25177 38795 25211
rect 38795 25177 38804 25211
rect 41420 25211 41472 25220
rect 38752 25168 38804 25177
rect 41420 25177 41429 25211
rect 41429 25177 41463 25211
rect 41463 25177 41472 25211
rect 42156 25245 42165 25279
rect 42165 25245 42199 25279
rect 42199 25245 42208 25279
rect 42156 25236 42208 25245
rect 45928 25279 45980 25288
rect 41420 25168 41472 25177
rect 41972 25168 42024 25220
rect 45928 25245 45937 25279
rect 45937 25245 45971 25279
rect 45971 25245 45980 25279
rect 45928 25236 45980 25245
rect 46112 25211 46164 25220
rect 46112 25177 46121 25211
rect 46121 25177 46155 25211
rect 46155 25177 46164 25211
rect 46112 25168 46164 25177
rect 28080 25100 28132 25152
rect 30380 25100 30432 25152
rect 31208 25100 31260 25152
rect 37096 25143 37148 25152
rect 37096 25109 37105 25143
rect 37105 25109 37139 25143
rect 37139 25109 37148 25143
rect 37096 25100 37148 25109
rect 37740 25143 37792 25152
rect 37740 25109 37749 25143
rect 37749 25109 37783 25143
rect 37783 25109 37792 25143
rect 37740 25100 37792 25109
rect 39120 25100 39172 25152
rect 42064 25100 42116 25152
rect 42892 25100 42944 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1768 24896 1820 24948
rect 23848 24896 23900 24948
rect 27896 24896 27948 24948
rect 29828 24939 29880 24948
rect 29828 24905 29837 24939
rect 29837 24905 29871 24939
rect 29871 24905 29880 24939
rect 29828 24896 29880 24905
rect 30932 24896 30984 24948
rect 30748 24828 30800 24880
rect 32496 24828 32548 24880
rect 34796 24828 34848 24880
rect 2964 24760 3016 24812
rect 3976 24760 4028 24812
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 22744 24760 22796 24812
rect 22928 24760 22980 24812
rect 27620 24803 27672 24812
rect 27620 24769 27629 24803
rect 27629 24769 27663 24803
rect 27663 24769 27672 24803
rect 27620 24760 27672 24769
rect 27804 24803 27856 24812
rect 27804 24769 27813 24803
rect 27813 24769 27847 24803
rect 27847 24769 27856 24803
rect 27804 24760 27856 24769
rect 27896 24803 27948 24812
rect 27896 24769 27905 24803
rect 27905 24769 27939 24803
rect 27939 24769 27948 24803
rect 28172 24803 28224 24812
rect 27896 24760 27948 24769
rect 28172 24769 28181 24803
rect 28181 24769 28215 24803
rect 28215 24769 28224 24803
rect 28172 24760 28224 24769
rect 30840 24760 30892 24812
rect 23112 24692 23164 24744
rect 23296 24624 23348 24676
rect 27436 24692 27488 24744
rect 30380 24692 30432 24744
rect 28080 24667 28132 24676
rect 28080 24633 28089 24667
rect 28089 24633 28123 24667
rect 28123 24633 28132 24667
rect 28080 24624 28132 24633
rect 30472 24624 30524 24676
rect 31024 24760 31076 24812
rect 31760 24760 31812 24812
rect 32956 24760 33008 24812
rect 35440 24803 35492 24812
rect 35440 24769 35449 24803
rect 35449 24769 35483 24803
rect 35483 24769 35492 24803
rect 35440 24760 35492 24769
rect 38752 24896 38804 24948
rect 39120 24896 39172 24948
rect 42156 24896 42208 24948
rect 38752 24803 38804 24812
rect 38752 24769 38786 24803
rect 38786 24769 38804 24803
rect 38752 24760 38804 24769
rect 35716 24735 35768 24744
rect 35716 24701 35725 24735
rect 35725 24701 35759 24735
rect 35759 24701 35768 24735
rect 35716 24692 35768 24701
rect 37188 24692 37240 24744
rect 38016 24692 38068 24744
rect 41144 24735 41196 24744
rect 41144 24701 41153 24735
rect 41153 24701 41187 24735
rect 41187 24701 41196 24735
rect 41144 24692 41196 24701
rect 41328 24760 41380 24812
rect 43260 24828 43312 24880
rect 42708 24760 42760 24812
rect 42892 24803 42944 24812
rect 42892 24769 42926 24803
rect 42926 24769 42944 24803
rect 42892 24760 42944 24769
rect 46020 24803 46072 24812
rect 46020 24769 46029 24803
rect 46029 24769 46063 24803
rect 46063 24769 46072 24803
rect 46020 24760 46072 24769
rect 47124 24803 47176 24812
rect 47124 24769 47133 24803
rect 47133 24769 47167 24803
rect 47167 24769 47176 24803
rect 47124 24760 47176 24769
rect 47400 24760 47452 24812
rect 47768 24760 47820 24812
rect 46848 24692 46900 24744
rect 35348 24556 35400 24608
rect 36084 24556 36136 24608
rect 41328 24556 41380 24608
rect 41972 24599 42024 24608
rect 41972 24565 41981 24599
rect 41981 24565 42015 24599
rect 42015 24565 42024 24599
rect 41972 24556 42024 24565
rect 45560 24624 45612 24676
rect 43904 24556 43956 24608
rect 45652 24556 45704 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 24952 24395 25004 24404
rect 24952 24361 24961 24395
rect 24961 24361 24995 24395
rect 24995 24361 25004 24395
rect 24952 24352 25004 24361
rect 27804 24352 27856 24404
rect 30380 24352 30432 24404
rect 23296 24259 23348 24268
rect 23296 24225 23305 24259
rect 23305 24225 23339 24259
rect 23339 24225 23348 24259
rect 23296 24216 23348 24225
rect 27712 24284 27764 24336
rect 31576 24352 31628 24404
rect 35440 24352 35492 24404
rect 35716 24352 35768 24404
rect 2044 24148 2096 24200
rect 22192 24148 22244 24200
rect 23020 24148 23072 24200
rect 23112 24080 23164 24132
rect 26148 24148 26200 24200
rect 27252 24191 27304 24200
rect 27252 24157 27262 24191
rect 27262 24157 27296 24191
rect 27296 24157 27304 24191
rect 27252 24148 27304 24157
rect 27436 24191 27488 24200
rect 27436 24157 27445 24191
rect 27445 24157 27479 24191
rect 27479 24157 27488 24191
rect 27436 24148 27488 24157
rect 27620 24191 27672 24200
rect 27620 24157 27634 24191
rect 27634 24157 27668 24191
rect 27668 24157 27672 24191
rect 28540 24191 28592 24200
rect 27620 24148 27672 24157
rect 26884 24080 26936 24132
rect 27528 24123 27580 24132
rect 27528 24089 27537 24123
rect 27537 24089 27571 24123
rect 27571 24089 27580 24123
rect 27528 24080 27580 24089
rect 28540 24157 28549 24191
rect 28549 24157 28583 24191
rect 28583 24157 28592 24191
rect 28540 24148 28592 24157
rect 28632 24191 28684 24200
rect 28632 24157 28641 24191
rect 28641 24157 28675 24191
rect 28675 24157 28684 24191
rect 28632 24148 28684 24157
rect 32956 24259 33008 24268
rect 32956 24225 32965 24259
rect 32965 24225 32999 24259
rect 32999 24225 33008 24259
rect 32956 24216 33008 24225
rect 30472 24148 30524 24200
rect 31760 24148 31812 24200
rect 34796 24148 34848 24200
rect 35348 24148 35400 24200
rect 37740 24284 37792 24336
rect 38752 24352 38804 24404
rect 41972 24352 42024 24404
rect 37924 24284 37976 24336
rect 41144 24284 41196 24336
rect 30380 24080 30432 24132
rect 33784 24080 33836 24132
rect 35992 24080 36044 24132
rect 37096 24148 37148 24200
rect 38660 24216 38712 24268
rect 39028 24259 39080 24268
rect 39028 24225 39037 24259
rect 39037 24225 39071 24259
rect 39071 24225 39080 24259
rect 39028 24216 39080 24225
rect 40132 24216 40184 24268
rect 42064 24216 42116 24268
rect 44180 24352 44232 24404
rect 46112 24352 46164 24404
rect 43260 24259 43312 24268
rect 43260 24225 43269 24259
rect 43269 24225 43303 24259
rect 43303 24225 43312 24259
rect 43260 24216 43312 24225
rect 37740 24191 37792 24200
rect 37740 24157 37749 24191
rect 37749 24157 37783 24191
rect 37783 24157 37792 24191
rect 37740 24148 37792 24157
rect 38844 24191 38896 24200
rect 23940 24055 23992 24064
rect 23940 24021 23949 24055
rect 23949 24021 23983 24055
rect 23983 24021 23992 24055
rect 23940 24012 23992 24021
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 25504 24012 25556 24064
rect 27804 24055 27856 24064
rect 27804 24021 27813 24055
rect 27813 24021 27847 24055
rect 27847 24021 27856 24055
rect 27804 24012 27856 24021
rect 30472 24012 30524 24064
rect 34612 24012 34664 24064
rect 35716 24012 35768 24064
rect 36912 24012 36964 24064
rect 37280 24055 37332 24064
rect 37280 24021 37289 24055
rect 37289 24021 37323 24055
rect 37323 24021 37332 24055
rect 37280 24012 37332 24021
rect 38844 24157 38853 24191
rect 38853 24157 38887 24191
rect 38887 24157 38896 24191
rect 38844 24148 38896 24157
rect 39120 24191 39172 24200
rect 39120 24157 39129 24191
rect 39129 24157 39163 24191
rect 39163 24157 39172 24191
rect 39120 24148 39172 24157
rect 42248 24191 42300 24200
rect 42248 24157 42257 24191
rect 42257 24157 42291 24191
rect 42291 24157 42300 24191
rect 42248 24148 42300 24157
rect 45652 24148 45704 24200
rect 46664 24148 46716 24200
rect 41144 24012 41196 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3516 23740 3568 23792
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 2228 23647 2280 23656
rect 2228 23613 2237 23647
rect 2237 23613 2271 23647
rect 2271 23613 2280 23647
rect 2228 23604 2280 23613
rect 2780 23647 2832 23656
rect 2780 23613 2789 23647
rect 2789 23613 2823 23647
rect 2823 23613 2832 23647
rect 2780 23604 2832 23613
rect 27252 23808 27304 23860
rect 27988 23808 28040 23860
rect 30380 23851 30432 23860
rect 30380 23817 30389 23851
rect 30389 23817 30423 23851
rect 30423 23817 30432 23851
rect 30380 23808 30432 23817
rect 30564 23808 30616 23860
rect 31300 23851 31352 23860
rect 31300 23817 31309 23851
rect 31309 23817 31343 23851
rect 31343 23817 31352 23851
rect 31300 23808 31352 23817
rect 33784 23851 33836 23860
rect 33784 23817 33793 23851
rect 33793 23817 33827 23851
rect 33827 23817 33836 23851
rect 33784 23808 33836 23817
rect 37740 23808 37792 23860
rect 40132 23851 40184 23860
rect 40132 23817 40157 23851
rect 40157 23817 40184 23851
rect 40132 23808 40184 23817
rect 40776 23808 40828 23860
rect 41328 23808 41380 23860
rect 22744 23740 22796 23792
rect 22376 23672 22428 23724
rect 30748 23740 30800 23792
rect 30932 23783 30984 23792
rect 30932 23749 30941 23783
rect 30941 23749 30975 23783
rect 30975 23749 30984 23783
rect 30932 23740 30984 23749
rect 35348 23740 35400 23792
rect 39948 23783 40000 23792
rect 39948 23749 39957 23783
rect 39957 23749 39991 23783
rect 39991 23749 40000 23783
rect 39948 23740 40000 23749
rect 44088 23740 44140 23792
rect 48044 23740 48096 23792
rect 24584 23672 24636 23724
rect 24860 23672 24912 23724
rect 25320 23715 25372 23724
rect 25320 23681 25329 23715
rect 25329 23681 25363 23715
rect 25363 23681 25372 23715
rect 25504 23715 25556 23724
rect 25320 23672 25372 23681
rect 25504 23681 25513 23715
rect 25513 23681 25547 23715
rect 25547 23681 25556 23715
rect 25504 23672 25556 23681
rect 26148 23715 26200 23724
rect 26148 23681 26157 23715
rect 26157 23681 26191 23715
rect 26191 23681 26200 23715
rect 26148 23672 26200 23681
rect 30472 23715 30524 23724
rect 22192 23647 22244 23656
rect 22192 23613 22201 23647
rect 22201 23613 22235 23647
rect 22235 23613 22244 23647
rect 22192 23604 22244 23613
rect 23204 23604 23256 23656
rect 26976 23604 27028 23656
rect 27712 23647 27764 23656
rect 27712 23613 27721 23647
rect 27721 23613 27755 23647
rect 27755 23613 27764 23647
rect 27712 23604 27764 23613
rect 28448 23604 28500 23656
rect 30472 23681 30481 23715
rect 30481 23681 30515 23715
rect 30515 23681 30524 23715
rect 30472 23672 30524 23681
rect 33692 23715 33744 23724
rect 33692 23681 33701 23715
rect 33701 23681 33735 23715
rect 33735 23681 33744 23715
rect 33692 23672 33744 23681
rect 34612 23672 34664 23724
rect 35992 23715 36044 23724
rect 35992 23681 36001 23715
rect 36001 23681 36035 23715
rect 36035 23681 36044 23715
rect 35992 23672 36044 23681
rect 36268 23715 36320 23724
rect 36268 23681 36277 23715
rect 36277 23681 36311 23715
rect 36311 23681 36320 23715
rect 36268 23672 36320 23681
rect 36360 23715 36412 23724
rect 36360 23681 36369 23715
rect 36369 23681 36403 23715
rect 36403 23681 36412 23715
rect 36360 23672 36412 23681
rect 37648 23672 37700 23724
rect 31208 23604 31260 23656
rect 37924 23604 37976 23656
rect 40040 23672 40092 23724
rect 41512 23715 41564 23724
rect 41512 23681 41522 23715
rect 41522 23681 41556 23715
rect 41556 23681 41564 23715
rect 41512 23672 41564 23681
rect 41696 23715 41748 23724
rect 41696 23681 41705 23715
rect 41705 23681 41739 23715
rect 41739 23681 41748 23715
rect 41696 23672 41748 23681
rect 42800 23672 42852 23724
rect 43904 23672 43956 23724
rect 42064 23604 42116 23656
rect 45376 23647 45428 23656
rect 45376 23613 45385 23647
rect 45385 23613 45419 23647
rect 45419 23613 45428 23647
rect 45376 23604 45428 23613
rect 45560 23647 45612 23656
rect 45560 23613 45569 23647
rect 45569 23613 45603 23647
rect 45603 23613 45612 23647
rect 45560 23604 45612 23613
rect 39488 23536 39540 23588
rect 41512 23536 41564 23588
rect 41972 23536 42024 23588
rect 23112 23511 23164 23520
rect 23112 23477 23121 23511
rect 23121 23477 23155 23511
rect 23155 23477 23164 23511
rect 23112 23468 23164 23477
rect 24952 23468 25004 23520
rect 28080 23468 28132 23520
rect 31392 23468 31444 23520
rect 36636 23468 36688 23520
rect 37556 23511 37608 23520
rect 37556 23477 37565 23511
rect 37565 23477 37599 23511
rect 37599 23477 37608 23511
rect 37556 23468 37608 23477
rect 38292 23468 38344 23520
rect 39120 23468 39172 23520
rect 40224 23468 40276 23520
rect 43812 23468 43864 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2228 23264 2280 23316
rect 24860 23264 24912 23316
rect 26148 23264 26200 23316
rect 27896 23264 27948 23316
rect 28540 23307 28592 23316
rect 28540 23273 28549 23307
rect 28549 23273 28583 23307
rect 28583 23273 28592 23307
rect 28540 23264 28592 23273
rect 34704 23264 34756 23316
rect 45560 23264 45612 23316
rect 23940 23128 23992 23180
rect 2412 23103 2464 23112
rect 2412 23069 2421 23103
rect 2421 23069 2455 23103
rect 2455 23069 2464 23103
rect 2412 23060 2464 23069
rect 23204 23103 23256 23112
rect 23204 23069 23213 23103
rect 23213 23069 23247 23103
rect 23247 23069 23256 23103
rect 23204 23060 23256 23069
rect 24400 23060 24452 23112
rect 24952 23103 25004 23112
rect 24952 23069 24986 23103
rect 24986 23069 25004 23103
rect 24952 23060 25004 23069
rect 26976 23103 27028 23112
rect 26976 23069 26985 23103
rect 26985 23069 27019 23103
rect 27019 23069 27028 23103
rect 26976 23060 27028 23069
rect 27068 23103 27120 23112
rect 27068 23069 27077 23103
rect 27077 23069 27111 23103
rect 27111 23069 27120 23103
rect 27068 23060 27120 23069
rect 27804 23196 27856 23248
rect 30564 23196 30616 23248
rect 27712 23128 27764 23180
rect 28632 23171 28684 23180
rect 28632 23137 28641 23171
rect 28641 23137 28675 23171
rect 28675 23137 28684 23171
rect 28632 23128 28684 23137
rect 31300 23196 31352 23248
rect 34796 23196 34848 23248
rect 37648 23196 37700 23248
rect 27804 23060 27856 23112
rect 28172 23103 28224 23112
rect 28172 23069 28178 23103
rect 28178 23069 28212 23103
rect 28212 23069 28224 23103
rect 28172 23060 28224 23069
rect 30656 23103 30708 23112
rect 30656 23069 30665 23103
rect 30665 23069 30699 23103
rect 30699 23069 30708 23103
rect 31300 23103 31352 23112
rect 30656 23060 30708 23069
rect 31300 23069 31309 23103
rect 31309 23069 31343 23103
rect 31343 23069 31352 23103
rect 31300 23060 31352 23069
rect 33692 23060 33744 23112
rect 33968 23060 34020 23112
rect 36636 23103 36688 23112
rect 36636 23069 36645 23103
rect 36645 23069 36679 23103
rect 36679 23069 36688 23103
rect 36636 23060 36688 23069
rect 36912 23103 36964 23112
rect 36912 23069 36921 23103
rect 36921 23069 36955 23103
rect 36955 23069 36964 23103
rect 36912 23060 36964 23069
rect 37556 23103 37608 23112
rect 37556 23069 37565 23103
rect 37565 23069 37599 23103
rect 37599 23069 37608 23103
rect 37556 23060 37608 23069
rect 38292 23103 38344 23112
rect 38292 23069 38301 23103
rect 38301 23069 38335 23103
rect 38335 23069 38344 23103
rect 38292 23060 38344 23069
rect 38476 23103 38528 23112
rect 38476 23069 38485 23103
rect 38485 23069 38519 23103
rect 38519 23069 38528 23103
rect 38476 23060 38528 23069
rect 27804 22924 27856 22976
rect 29920 22924 29972 22976
rect 34612 22992 34664 23044
rect 35348 22992 35400 23044
rect 37280 22992 37332 23044
rect 39304 22992 39356 23044
rect 39948 22992 40000 23044
rect 41696 23128 41748 23180
rect 42708 23128 42760 23180
rect 43260 23171 43312 23180
rect 43260 23137 43269 23171
rect 43269 23137 43303 23171
rect 43303 23137 43312 23171
rect 43260 23128 43312 23137
rect 44088 23171 44140 23180
rect 44088 23137 44097 23171
rect 44097 23137 44131 23171
rect 44131 23137 44140 23171
rect 44088 23128 44140 23137
rect 44180 23171 44232 23180
rect 44180 23137 44189 23171
rect 44189 23137 44223 23171
rect 44223 23137 44232 23171
rect 44180 23128 44232 23137
rect 40132 23060 40184 23112
rect 40776 23103 40828 23112
rect 40776 23069 40785 23103
rect 40785 23069 40819 23103
rect 40819 23069 40828 23103
rect 40776 23060 40828 23069
rect 41052 23103 41104 23112
rect 41052 23069 41061 23103
rect 41061 23069 41095 23103
rect 41095 23069 41104 23103
rect 41052 23060 41104 23069
rect 41604 23103 41656 23112
rect 41604 23069 41613 23103
rect 41613 23069 41647 23103
rect 41647 23069 41656 23103
rect 41604 23060 41656 23069
rect 43812 23103 43864 23112
rect 43812 23069 43821 23103
rect 43821 23069 43855 23103
rect 43855 23069 43864 23103
rect 43812 23060 43864 23069
rect 43904 23060 43956 23112
rect 45652 23103 45704 23112
rect 40224 23035 40276 23044
rect 40224 23001 40233 23035
rect 40233 23001 40267 23035
rect 40267 23001 40276 23035
rect 40224 22992 40276 23001
rect 41236 22992 41288 23044
rect 44272 22992 44324 23044
rect 31116 22924 31168 22976
rect 37372 22967 37424 22976
rect 37372 22933 37381 22967
rect 37381 22933 37415 22967
rect 37415 22933 37424 22967
rect 37372 22924 37424 22933
rect 37464 22924 37516 22976
rect 38384 22967 38436 22976
rect 38384 22933 38393 22967
rect 38393 22933 38427 22967
rect 38427 22933 38436 22967
rect 38384 22924 38436 22933
rect 40776 22967 40828 22976
rect 40776 22933 40785 22967
rect 40785 22933 40819 22967
rect 40819 22933 40828 22967
rect 40776 22924 40828 22933
rect 44088 22924 44140 22976
rect 45652 23069 45661 23103
rect 45661 23069 45695 23103
rect 45695 23069 45704 23103
rect 45652 23060 45704 23069
rect 46480 23103 46532 23112
rect 46480 23069 46489 23103
rect 46489 23069 46523 23103
rect 46523 23069 46532 23103
rect 46480 23060 46532 23069
rect 47124 22992 47176 23044
rect 48320 23035 48372 23044
rect 48320 23001 48329 23035
rect 48329 23001 48363 23035
rect 48363 23001 48372 23035
rect 48320 22992 48372 23001
rect 44456 22924 44508 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 27068 22720 27120 22772
rect 2412 22652 2464 22704
rect 5448 22652 5500 22704
rect 23204 22627 23256 22636
rect 23204 22593 23213 22627
rect 23213 22593 23247 22627
rect 23247 22593 23256 22627
rect 23204 22584 23256 22593
rect 23296 22584 23348 22636
rect 26424 22627 26476 22636
rect 26424 22593 26433 22627
rect 26433 22593 26467 22627
rect 26467 22593 26476 22627
rect 26424 22584 26476 22593
rect 27620 22720 27672 22772
rect 28448 22763 28500 22772
rect 28448 22729 28457 22763
rect 28457 22729 28491 22763
rect 28491 22729 28500 22763
rect 28448 22720 28500 22729
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 28172 22584 28224 22636
rect 30472 22652 30524 22704
rect 30380 22627 30432 22636
rect 27528 22448 27580 22500
rect 27804 22491 27856 22500
rect 27804 22457 27813 22491
rect 27813 22457 27847 22491
rect 27847 22457 27856 22491
rect 27804 22448 27856 22457
rect 30380 22593 30389 22627
rect 30389 22593 30423 22627
rect 30423 22593 30432 22627
rect 30380 22584 30432 22593
rect 30748 22652 30800 22704
rect 37464 22720 37516 22772
rect 37556 22720 37608 22772
rect 36636 22652 36688 22704
rect 37372 22652 37424 22704
rect 29920 22559 29972 22568
rect 29920 22525 29929 22559
rect 29929 22525 29963 22559
rect 29963 22525 29972 22559
rect 30932 22584 30984 22636
rect 31392 22627 31444 22636
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 31484 22627 31536 22636
rect 31484 22593 31493 22627
rect 31493 22593 31527 22627
rect 31527 22593 31536 22627
rect 31484 22584 31536 22593
rect 33140 22584 33192 22636
rect 33876 22627 33928 22636
rect 33876 22593 33910 22627
rect 33910 22593 33928 22627
rect 36360 22627 36412 22636
rect 33876 22584 33928 22593
rect 29920 22516 29972 22525
rect 31116 22516 31168 22568
rect 30656 22448 30708 22500
rect 23388 22380 23440 22432
rect 29460 22423 29512 22432
rect 29460 22389 29469 22423
rect 29469 22389 29503 22423
rect 29503 22389 29512 22423
rect 29460 22380 29512 22389
rect 30472 22380 30524 22432
rect 32496 22380 32548 22432
rect 34704 22380 34756 22432
rect 36360 22593 36369 22627
rect 36369 22593 36403 22627
rect 36403 22593 36412 22627
rect 36360 22584 36412 22593
rect 36268 22516 36320 22568
rect 36544 22584 36596 22636
rect 37740 22627 37792 22636
rect 37740 22593 37749 22627
rect 37749 22593 37783 22627
rect 37783 22593 37792 22627
rect 37740 22584 37792 22593
rect 36820 22516 36872 22568
rect 38844 22584 38896 22636
rect 40040 22720 40092 22772
rect 41696 22720 41748 22772
rect 44088 22720 44140 22772
rect 47124 22763 47176 22772
rect 47124 22729 47133 22763
rect 47133 22729 47167 22763
rect 47167 22729 47176 22763
rect 47124 22720 47176 22729
rect 39120 22627 39172 22636
rect 39120 22593 39129 22627
rect 39129 22593 39163 22627
rect 39163 22593 39172 22627
rect 39120 22584 39172 22593
rect 39304 22627 39356 22636
rect 39304 22593 39313 22627
rect 39313 22593 39347 22627
rect 39347 22593 39356 22627
rect 39304 22584 39356 22593
rect 39488 22627 39540 22636
rect 39488 22593 39497 22627
rect 39497 22593 39531 22627
rect 39531 22593 39540 22627
rect 39488 22584 39540 22593
rect 41604 22652 41656 22704
rect 44180 22695 44232 22704
rect 44180 22661 44189 22695
rect 44189 22661 44223 22695
rect 44223 22661 44232 22695
rect 44180 22652 44232 22661
rect 45376 22652 45428 22704
rect 46480 22652 46532 22704
rect 40776 22584 40828 22636
rect 43352 22627 43404 22636
rect 43352 22593 43361 22627
rect 43361 22593 43395 22627
rect 43395 22593 43404 22627
rect 43352 22584 43404 22593
rect 44456 22627 44508 22636
rect 44456 22593 44465 22627
rect 44465 22593 44499 22627
rect 44499 22593 44508 22627
rect 44456 22584 44508 22593
rect 45100 22627 45152 22636
rect 45100 22593 45109 22627
rect 45109 22593 45143 22627
rect 45143 22593 45152 22627
rect 45100 22584 45152 22593
rect 47032 22627 47084 22636
rect 47032 22593 47041 22627
rect 47041 22593 47075 22627
rect 47075 22593 47084 22627
rect 47032 22584 47084 22593
rect 39028 22516 39080 22568
rect 44272 22516 44324 22568
rect 37740 22448 37792 22500
rect 43996 22448 44048 22500
rect 41512 22380 41564 22432
rect 45652 22380 45704 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 26976 22176 27028 22228
rect 30380 22176 30432 22228
rect 31116 22219 31168 22228
rect 31116 22185 31125 22219
rect 31125 22185 31159 22219
rect 31159 22185 31168 22219
rect 31116 22176 31168 22185
rect 33876 22176 33928 22228
rect 36636 22176 36688 22228
rect 41512 22176 41564 22228
rect 41604 22176 41656 22228
rect 42708 22176 42760 22228
rect 2780 22083 2832 22092
rect 2780 22049 2789 22083
rect 2789 22049 2823 22083
rect 2823 22049 2832 22083
rect 2780 22040 2832 22049
rect 26240 22040 26292 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 22836 21972 22888 22024
rect 23204 21972 23256 22024
rect 29736 22015 29788 22024
rect 1768 21947 1820 21956
rect 1768 21913 1777 21947
rect 1777 21913 1811 21947
rect 1811 21913 1820 21947
rect 1768 21904 1820 21913
rect 29736 21981 29745 22015
rect 29745 21981 29779 22015
rect 29779 21981 29788 22015
rect 29736 21972 29788 21981
rect 34796 22040 34848 22092
rect 34704 21972 34756 22024
rect 35348 21972 35400 22024
rect 37280 22015 37332 22024
rect 37280 21981 37289 22015
rect 37289 21981 37323 22015
rect 37323 21981 37332 22015
rect 37280 21972 37332 21981
rect 40500 21972 40552 22024
rect 41144 22015 41196 22024
rect 41144 21981 41153 22015
rect 41153 21981 41187 22015
rect 41187 21981 41196 22015
rect 41604 22015 41656 22024
rect 41144 21972 41196 21981
rect 29460 21904 29512 21956
rect 33968 21904 34020 21956
rect 34336 21947 34388 21956
rect 34336 21913 34345 21947
rect 34345 21913 34379 21947
rect 34379 21913 34388 21947
rect 34336 21904 34388 21913
rect 34612 21904 34664 21956
rect 38384 21904 38436 21956
rect 41604 21981 41613 22015
rect 41613 21981 41647 22015
rect 41647 21981 41656 22015
rect 41604 21972 41656 21981
rect 43352 22176 43404 22228
rect 43996 22083 44048 22092
rect 43996 22049 44005 22083
rect 44005 22049 44039 22083
rect 44039 22049 44048 22083
rect 43996 22040 44048 22049
rect 44088 21972 44140 22024
rect 46480 22015 46532 22024
rect 46480 21981 46489 22015
rect 46489 21981 46523 22015
rect 46523 21981 46532 22015
rect 46480 21972 46532 21981
rect 42064 21904 42116 21956
rect 47124 21904 47176 21956
rect 48320 21947 48372 21956
rect 48320 21913 48329 21947
rect 48329 21913 48363 21947
rect 48363 21913 48372 21947
rect 48320 21904 48372 21913
rect 23204 21836 23256 21888
rect 23388 21836 23440 21888
rect 37740 21836 37792 21888
rect 41788 21836 41840 21888
rect 44180 21836 44232 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1768 21632 1820 21684
rect 22836 21675 22888 21684
rect 22836 21641 22845 21675
rect 22845 21641 22879 21675
rect 22879 21641 22888 21675
rect 22836 21632 22888 21641
rect 23480 21632 23532 21684
rect 26424 21632 26476 21684
rect 30196 21632 30248 21684
rect 31392 21632 31444 21684
rect 38476 21632 38528 21684
rect 1584 21496 1636 21548
rect 2964 21496 3016 21548
rect 30472 21564 30524 21616
rect 47124 21675 47176 21684
rect 47124 21641 47133 21675
rect 47133 21641 47167 21675
rect 47167 21641 47176 21675
rect 47124 21632 47176 21641
rect 42064 21607 42116 21616
rect 42064 21573 42073 21607
rect 42073 21573 42107 21607
rect 42107 21573 42116 21607
rect 42064 21564 42116 21573
rect 46480 21564 46532 21616
rect 23112 21496 23164 21548
rect 23480 21496 23532 21548
rect 23756 21539 23808 21548
rect 23756 21505 23765 21539
rect 23765 21505 23799 21539
rect 23799 21505 23808 21539
rect 23756 21496 23808 21505
rect 24032 21496 24084 21548
rect 24400 21539 24452 21548
rect 24400 21505 24409 21539
rect 24409 21505 24443 21539
rect 24443 21505 24452 21539
rect 24400 21496 24452 21505
rect 26884 21496 26936 21548
rect 28264 21496 28316 21548
rect 31484 21496 31536 21548
rect 37648 21539 37700 21548
rect 37648 21505 37657 21539
rect 37657 21505 37691 21539
rect 37691 21505 37700 21539
rect 37648 21496 37700 21505
rect 41696 21539 41748 21548
rect 41696 21505 41705 21539
rect 41705 21505 41739 21539
rect 41739 21505 41748 21539
rect 41696 21496 41748 21505
rect 41788 21496 41840 21548
rect 44272 21496 44324 21548
rect 47032 21539 47084 21548
rect 47032 21505 47041 21539
rect 47041 21505 47075 21539
rect 47075 21505 47084 21539
rect 47032 21496 47084 21505
rect 2320 21360 2372 21412
rect 2688 21360 2740 21412
rect 23848 21360 23900 21412
rect 37740 21428 37792 21480
rect 41420 21428 41472 21480
rect 44180 21471 44232 21480
rect 44180 21437 44189 21471
rect 44189 21437 44223 21471
rect 44223 21437 44232 21471
rect 44180 21428 44232 21437
rect 27436 21292 27488 21344
rect 29920 21292 29972 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 23756 21088 23808 21140
rect 28264 21131 28316 21140
rect 28264 21097 28273 21131
rect 28273 21097 28307 21131
rect 28307 21097 28316 21131
rect 28264 21088 28316 21097
rect 31392 21088 31444 21140
rect 31484 21088 31536 21140
rect 44640 21131 44692 21140
rect 44640 21097 44649 21131
rect 44649 21097 44683 21131
rect 44683 21097 44692 21131
rect 44640 21088 44692 21097
rect 45100 21088 45152 21140
rect 23112 21020 23164 21072
rect 23204 20995 23256 21004
rect 23204 20961 23213 20995
rect 23213 20961 23247 20995
rect 23247 20961 23256 20995
rect 23204 20952 23256 20961
rect 24400 21020 24452 21072
rect 2044 20884 2096 20936
rect 23388 20884 23440 20936
rect 42708 20952 42760 21004
rect 29736 20927 29788 20936
rect 23848 20816 23900 20868
rect 25320 20816 25372 20868
rect 26700 20816 26752 20868
rect 26332 20748 26384 20800
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 31300 20884 31352 20936
rect 32312 20884 32364 20936
rect 33048 20884 33100 20936
rect 27528 20816 27580 20868
rect 29828 20816 29880 20868
rect 31852 20859 31904 20868
rect 31852 20825 31886 20859
rect 31886 20825 31904 20859
rect 31852 20816 31904 20825
rect 35348 20816 35400 20868
rect 42984 20816 43036 20868
rect 28172 20748 28224 20800
rect 36268 20791 36320 20800
rect 36268 20757 36277 20791
rect 36277 20757 36311 20791
rect 36311 20757 36320 20791
rect 36268 20748 36320 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 23296 20587 23348 20596
rect 23296 20553 23305 20587
rect 23305 20553 23339 20587
rect 23339 20553 23348 20587
rect 23296 20544 23348 20553
rect 26700 20544 26752 20596
rect 28172 20587 28224 20596
rect 28172 20553 28181 20587
rect 28181 20553 28215 20587
rect 28215 20553 28224 20587
rect 28172 20544 28224 20553
rect 29828 20544 29880 20596
rect 31852 20544 31904 20596
rect 35348 20587 35400 20596
rect 35348 20553 35357 20587
rect 35357 20553 35391 20587
rect 35391 20553 35400 20587
rect 35348 20544 35400 20553
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 23112 20408 23164 20460
rect 23480 20408 23532 20460
rect 26240 20451 26292 20460
rect 26240 20417 26249 20451
rect 26249 20417 26283 20451
rect 26283 20417 26292 20451
rect 26240 20408 26292 20417
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 28264 20408 28316 20460
rect 29920 20451 29972 20460
rect 29920 20417 29929 20451
rect 29929 20417 29963 20451
rect 29963 20417 29972 20451
rect 29920 20408 29972 20417
rect 30196 20451 30248 20460
rect 30196 20417 30205 20451
rect 30205 20417 30239 20451
rect 30239 20417 30248 20451
rect 30196 20408 30248 20417
rect 31484 20408 31536 20460
rect 34336 20476 34388 20528
rect 38476 20544 38528 20596
rect 42984 20587 43036 20596
rect 32312 20451 32364 20460
rect 32312 20417 32321 20451
rect 32321 20417 32355 20451
rect 32355 20417 32364 20451
rect 32312 20408 32364 20417
rect 32864 20408 32916 20460
rect 33876 20408 33928 20460
rect 34612 20451 34664 20460
rect 34612 20417 34621 20451
rect 34621 20417 34655 20451
rect 34655 20417 34664 20451
rect 34612 20408 34664 20417
rect 34796 20451 34848 20460
rect 34796 20417 34805 20451
rect 34805 20417 34839 20451
rect 34839 20417 34848 20451
rect 34796 20408 34848 20417
rect 38200 20476 38252 20528
rect 35808 20451 35860 20460
rect 2504 20340 2556 20392
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 26332 20383 26384 20392
rect 26332 20349 26341 20383
rect 26341 20349 26375 20383
rect 26375 20349 26384 20383
rect 26332 20340 26384 20349
rect 26976 20340 27028 20392
rect 35808 20417 35817 20451
rect 35817 20417 35851 20451
rect 35851 20417 35860 20451
rect 35808 20408 35860 20417
rect 36084 20408 36136 20460
rect 36360 20408 36412 20460
rect 36268 20340 36320 20392
rect 37280 20408 37332 20460
rect 38016 20451 38068 20460
rect 38016 20417 38050 20451
rect 38050 20417 38068 20451
rect 41604 20476 41656 20528
rect 42984 20553 42993 20587
rect 42993 20553 43027 20587
rect 43027 20553 43036 20587
rect 42984 20544 43036 20553
rect 38016 20408 38068 20417
rect 41328 20408 41380 20460
rect 27528 20247 27580 20256
rect 27528 20213 27537 20247
rect 27537 20213 27571 20247
rect 27571 20213 27580 20247
rect 27528 20204 27580 20213
rect 33048 20204 33100 20256
rect 33692 20247 33744 20256
rect 33692 20213 33701 20247
rect 33701 20213 33735 20247
rect 33735 20213 33744 20247
rect 33692 20204 33744 20213
rect 34244 20204 34296 20256
rect 35992 20204 36044 20256
rect 36544 20247 36596 20256
rect 36544 20213 36553 20247
rect 36553 20213 36587 20247
rect 36587 20213 36596 20247
rect 36544 20204 36596 20213
rect 37740 20204 37792 20256
rect 38108 20204 38160 20256
rect 40500 20272 40552 20324
rect 39120 20247 39172 20256
rect 39120 20213 39129 20247
rect 39129 20213 39163 20247
rect 39163 20213 39172 20247
rect 39120 20204 39172 20213
rect 41880 20247 41932 20256
rect 41880 20213 41889 20247
rect 41889 20213 41923 20247
rect 41923 20213 41932 20247
rect 41880 20204 41932 20213
rect 43444 20451 43496 20460
rect 43444 20417 43453 20451
rect 43453 20417 43487 20451
rect 43487 20417 43496 20451
rect 43444 20408 43496 20417
rect 44088 20451 44140 20460
rect 44088 20417 44097 20451
rect 44097 20417 44131 20451
rect 44131 20417 44140 20451
rect 44088 20408 44140 20417
rect 43352 20272 43404 20324
rect 44640 20408 44692 20460
rect 47032 20451 47084 20460
rect 47032 20417 47041 20451
rect 47041 20417 47075 20451
rect 47075 20417 47084 20451
rect 47032 20408 47084 20417
rect 47308 20408 47360 20460
rect 43996 20204 44048 20256
rect 46664 20204 46716 20256
rect 47952 20247 48004 20256
rect 47952 20213 47961 20247
rect 47961 20213 47995 20247
rect 47995 20213 48004 20247
rect 47952 20204 48004 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2504 20043 2556 20052
rect 2504 20009 2513 20043
rect 2513 20009 2547 20043
rect 2547 20009 2556 20043
rect 2504 20000 2556 20009
rect 32864 20043 32916 20052
rect 32864 20009 32873 20043
rect 32873 20009 32907 20043
rect 32907 20009 32916 20043
rect 32864 20000 32916 20009
rect 33968 20000 34020 20052
rect 34796 20000 34848 20052
rect 35808 20000 35860 20052
rect 35900 20000 35952 20052
rect 36176 20000 36228 20052
rect 38016 20000 38068 20052
rect 39028 20043 39080 20052
rect 34244 19932 34296 19984
rect 2136 19796 2188 19848
rect 3240 19796 3292 19848
rect 33692 19864 33744 19916
rect 33324 19839 33376 19848
rect 33324 19805 33333 19839
rect 33333 19805 33367 19839
rect 33367 19805 33376 19839
rect 33324 19796 33376 19805
rect 34612 19796 34664 19848
rect 33876 19728 33928 19780
rect 34336 19728 34388 19780
rect 34704 19728 34756 19780
rect 35348 19839 35400 19848
rect 35348 19805 35357 19839
rect 35357 19805 35391 19839
rect 35391 19805 35400 19839
rect 35348 19796 35400 19805
rect 35900 19796 35952 19848
rect 36268 19907 36320 19916
rect 36268 19873 36277 19907
rect 36277 19873 36311 19907
rect 36311 19873 36320 19907
rect 36268 19864 36320 19873
rect 38200 19932 38252 19984
rect 39028 20009 39037 20043
rect 39037 20009 39071 20043
rect 39071 20009 39080 20043
rect 39028 20000 39080 20009
rect 41328 20043 41380 20052
rect 41328 20009 41337 20043
rect 41337 20009 41371 20043
rect 41371 20009 41380 20043
rect 41328 20000 41380 20009
rect 41972 20043 42024 20052
rect 41972 20009 41981 20043
rect 41981 20009 42015 20043
rect 42015 20009 42024 20043
rect 41972 20000 42024 20009
rect 43444 20000 43496 20052
rect 40132 19932 40184 19984
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 38476 19839 38528 19848
rect 38476 19805 38485 19839
rect 38485 19805 38519 19839
rect 38519 19805 38528 19839
rect 39120 19864 39172 19916
rect 38476 19796 38528 19805
rect 39488 19796 39540 19848
rect 40132 19796 40184 19848
rect 41236 19839 41288 19848
rect 41236 19805 41245 19839
rect 41245 19805 41279 19839
rect 41279 19805 41288 19839
rect 41236 19796 41288 19805
rect 41328 19839 41380 19848
rect 41328 19805 41337 19839
rect 41337 19805 41371 19839
rect 41371 19805 41380 19839
rect 41880 19839 41932 19848
rect 41328 19796 41380 19805
rect 41880 19805 41889 19839
rect 41889 19805 41923 19839
rect 41923 19805 41932 19839
rect 41880 19796 41932 19805
rect 43168 19839 43220 19848
rect 43168 19805 43177 19839
rect 43177 19805 43211 19839
rect 43211 19805 43220 19839
rect 43168 19796 43220 19805
rect 43352 19839 43404 19848
rect 43352 19805 43361 19839
rect 43361 19805 43395 19839
rect 43395 19805 43404 19839
rect 44640 19864 44692 19916
rect 47952 19932 48004 19984
rect 46664 19907 46716 19916
rect 46664 19873 46673 19907
rect 46673 19873 46707 19907
rect 46707 19873 46716 19907
rect 46664 19864 46716 19873
rect 48228 19907 48280 19916
rect 48228 19873 48237 19907
rect 48237 19873 48271 19907
rect 48271 19873 48280 19907
rect 48228 19864 48280 19873
rect 43352 19796 43404 19805
rect 44088 19796 44140 19848
rect 34796 19660 34848 19712
rect 34980 19660 35032 19712
rect 35808 19703 35860 19712
rect 35808 19669 35817 19703
rect 35817 19669 35851 19703
rect 35851 19669 35860 19703
rect 35808 19660 35860 19669
rect 36820 19703 36872 19712
rect 36820 19669 36829 19703
rect 36829 19669 36863 19703
rect 36863 19669 36872 19703
rect 36820 19660 36872 19669
rect 38200 19660 38252 19712
rect 40040 19703 40092 19712
rect 40040 19669 40049 19703
rect 40049 19669 40083 19703
rect 40083 19669 40092 19703
rect 40040 19660 40092 19669
rect 40592 19728 40644 19780
rect 41696 19660 41748 19712
rect 44364 19660 44416 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 33324 19456 33376 19508
rect 35164 19456 35216 19508
rect 35440 19456 35492 19508
rect 34980 19388 35032 19440
rect 33048 19363 33100 19372
rect 33048 19329 33057 19363
rect 33057 19329 33091 19363
rect 33091 19329 33100 19363
rect 33048 19320 33100 19329
rect 35716 19388 35768 19440
rect 36360 19456 36412 19508
rect 38108 19456 38160 19508
rect 38292 19456 38344 19508
rect 41236 19499 41288 19508
rect 35992 19388 36044 19440
rect 33508 19295 33560 19304
rect 33508 19261 33517 19295
rect 33517 19261 33551 19295
rect 33551 19261 33560 19295
rect 33508 19252 33560 19261
rect 33968 19295 34020 19304
rect 33968 19261 33977 19295
rect 33977 19261 34011 19295
rect 34011 19261 34020 19295
rect 33968 19252 34020 19261
rect 35808 19320 35860 19372
rect 35164 19295 35216 19304
rect 35164 19261 35173 19295
rect 35173 19261 35207 19295
rect 35207 19261 35216 19295
rect 35164 19252 35216 19261
rect 38752 19388 38804 19440
rect 39948 19388 40000 19440
rect 41236 19465 41245 19499
rect 41245 19465 41279 19499
rect 41279 19465 41288 19499
rect 41236 19456 41288 19465
rect 43168 19456 43220 19508
rect 43812 19456 43864 19508
rect 38936 19320 38988 19372
rect 38568 19252 38620 19304
rect 39120 19320 39172 19372
rect 39488 19363 39540 19372
rect 39488 19329 39497 19363
rect 39497 19329 39531 19363
rect 39531 19329 39540 19363
rect 39488 19320 39540 19329
rect 40040 19320 40092 19372
rect 40684 19320 40736 19372
rect 41880 19320 41932 19372
rect 40224 19252 40276 19304
rect 43812 19320 43864 19372
rect 44364 19363 44416 19372
rect 44364 19329 44373 19363
rect 44373 19329 44407 19363
rect 44407 19329 44416 19363
rect 44364 19320 44416 19329
rect 47216 19320 47268 19372
rect 47676 19320 47728 19372
rect 38660 19184 38712 19236
rect 39672 19159 39724 19168
rect 39672 19125 39681 19159
rect 39681 19125 39715 19159
rect 39715 19125 39724 19159
rect 39672 19116 39724 19125
rect 39948 19116 40000 19168
rect 44272 19252 44324 19304
rect 47124 19159 47176 19168
rect 47124 19125 47133 19159
rect 47133 19125 47167 19159
rect 47167 19125 47176 19159
rect 47124 19116 47176 19125
rect 47952 19159 48004 19168
rect 47952 19125 47961 19159
rect 47961 19125 47995 19159
rect 47995 19125 48004 19159
rect 47952 19116 48004 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 34336 18912 34388 18964
rect 35716 18955 35768 18964
rect 35716 18921 35725 18955
rect 35725 18921 35759 18955
rect 35759 18921 35768 18955
rect 35716 18912 35768 18921
rect 38936 18955 38988 18964
rect 38936 18921 38945 18955
rect 38945 18921 38979 18955
rect 38979 18921 38988 18955
rect 38936 18912 38988 18921
rect 43812 18955 43864 18964
rect 43812 18921 43821 18955
rect 43821 18921 43855 18955
rect 43855 18921 43864 18955
rect 43812 18912 43864 18921
rect 2044 18708 2096 18760
rect 35624 18776 35676 18828
rect 36176 18776 36228 18828
rect 39488 18844 39540 18896
rect 40592 18887 40644 18896
rect 40592 18853 40601 18887
rect 40601 18853 40635 18887
rect 40635 18853 40644 18887
rect 40592 18844 40644 18853
rect 34244 18708 34296 18760
rect 36544 18708 36596 18760
rect 39028 18776 39080 18828
rect 39672 18776 39724 18828
rect 38660 18708 38712 18760
rect 38752 18751 38804 18760
rect 38752 18717 38761 18751
rect 38761 18717 38795 18751
rect 38795 18717 38804 18751
rect 40224 18751 40276 18760
rect 38752 18708 38804 18717
rect 40224 18717 40233 18751
rect 40233 18717 40267 18751
rect 40267 18717 40276 18751
rect 40224 18708 40276 18717
rect 44364 18776 44416 18828
rect 47952 18844 48004 18896
rect 47124 18776 47176 18828
rect 48228 18819 48280 18828
rect 48228 18785 48237 18819
rect 48237 18785 48271 18819
rect 48271 18785 48280 18819
rect 48228 18776 48280 18785
rect 43996 18751 44048 18760
rect 43996 18717 44005 18751
rect 44005 18717 44039 18751
rect 44039 18717 44048 18751
rect 43996 18708 44048 18717
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 35440 18411 35492 18420
rect 35440 18377 35449 18411
rect 35449 18377 35483 18411
rect 35483 18377 35492 18411
rect 35440 18368 35492 18377
rect 38568 18411 38620 18420
rect 38568 18377 38577 18411
rect 38577 18377 38611 18411
rect 38611 18377 38620 18411
rect 38568 18368 38620 18377
rect 38660 18368 38712 18420
rect 40224 18368 40276 18420
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 36820 18232 36872 18284
rect 38752 18232 38804 18284
rect 41972 18232 42024 18284
rect 47492 18232 47544 18284
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 35624 18164 35676 18216
rect 40132 18207 40184 18216
rect 40132 18173 40141 18207
rect 40141 18173 40175 18207
rect 40175 18173 40184 18207
rect 40132 18164 40184 18173
rect 47860 18071 47912 18080
rect 47860 18037 47869 18071
rect 47869 18037 47903 18071
rect 47903 18037 47912 18071
rect 47860 18028 47912 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2228 17824 2280 17876
rect 47860 17688 47912 17740
rect 48228 17731 48280 17740
rect 48228 17697 48237 17731
rect 48237 17697 48271 17731
rect 48271 17697 48280 17731
rect 48228 17688 48280 17697
rect 2504 17620 2556 17672
rect 4620 17620 4672 17672
rect 46480 17663 46532 17672
rect 46480 17629 46489 17663
rect 46489 17629 46523 17663
rect 46523 17629 46532 17663
rect 46480 17620 46532 17629
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2872 17212 2924 17264
rect 46480 17144 46532 17196
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 46480 16940 46532 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2044 16736 2096 16788
rect 2596 16600 2648 16652
rect 3792 16600 3844 16652
rect 46480 16643 46532 16652
rect 46480 16609 46489 16643
rect 46489 16609 46523 16643
rect 46523 16609 46532 16643
rect 46480 16600 46532 16609
rect 48228 16643 48280 16652
rect 48228 16609 48237 16643
rect 48237 16609 48271 16643
rect 48271 16609 48280 16643
rect 48228 16600 48280 16609
rect 2872 16507 2924 16516
rect 2872 16473 2881 16507
rect 2881 16473 2915 16507
rect 2915 16473 2924 16507
rect 2872 16464 2924 16473
rect 47860 16464 47912 16516
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 47860 16235 47912 16244
rect 47860 16201 47869 16235
rect 47869 16201 47903 16235
rect 47903 16201 47912 16235
rect 47860 16192 47912 16201
rect 47768 16099 47820 16108
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 2136 15444 2188 15496
rect 2596 15444 2648 15496
rect 47676 15487 47728 15496
rect 47676 15453 47685 15487
rect 47685 15453 47719 15487
rect 47719 15453 47728 15487
rect 47676 15444 47728 15453
rect 2228 15308 2280 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2228 15079 2280 15088
rect 2228 15045 2237 15079
rect 2237 15045 2271 15079
rect 2271 15045 2280 15079
rect 2228 15036 2280 15045
rect 1952 14968 2004 15020
rect 47492 14968 47544 15020
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 46664 14764 46716 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 47676 14492 47728 14544
rect 46664 14467 46716 14476
rect 46664 14433 46673 14467
rect 46673 14433 46707 14467
rect 46707 14433 46716 14467
rect 46664 14424 46716 14433
rect 48228 14467 48280 14476
rect 48228 14433 48237 14467
rect 48237 14433 48271 14467
rect 48271 14433 48280 14467
rect 48228 14424 48280 14433
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 1768 14331 1820 14340
rect 1768 14297 1777 14331
rect 1777 14297 1811 14331
rect 1811 14297 1820 14331
rect 1768 14288 1820 14297
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1768 14016 1820 14068
rect 1584 13880 1636 13932
rect 2688 13880 2740 13932
rect 3056 13880 3108 13932
rect 47492 13880 47544 13932
rect 47124 13719 47176 13728
rect 47124 13685 47133 13719
rect 47133 13685 47167 13719
rect 47167 13685 47176 13719
rect 47124 13676 47176 13685
rect 47952 13719 48004 13728
rect 47952 13685 47961 13719
rect 47961 13685 47995 13719
rect 47995 13685 48004 13719
rect 47952 13676 48004 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 47952 13404 48004 13456
rect 47124 13336 47176 13388
rect 48228 13379 48280 13388
rect 48228 13345 48237 13379
rect 48237 13345 48271 13379
rect 48271 13345 48280 13379
rect 48228 13336 48280 13345
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 46940 12792 46992 12844
rect 47124 12631 47176 12640
rect 47124 12597 47133 12631
rect 47133 12597 47167 12631
rect 47167 12597 47176 12631
rect 47124 12588 47176 12597
rect 47952 12631 48004 12640
rect 47952 12597 47961 12631
rect 47961 12597 47995 12631
rect 47995 12597 48004 12631
rect 47952 12588 48004 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 47952 12316 48004 12368
rect 47124 12248 47176 12300
rect 48228 12291 48280 12300
rect 48228 12257 48237 12291
rect 48237 12257 48271 12291
rect 48271 12257 48280 12291
rect 48228 12248 48280 12257
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2320 11772 2372 11824
rect 47032 11747 47084 11756
rect 47032 11713 47041 11747
rect 47041 11713 47075 11747
rect 47075 11713 47084 11747
rect 47032 11704 47084 11713
rect 2320 11636 2372 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 46664 11500 46716 11552
rect 47952 11543 48004 11552
rect 47952 11509 47961 11543
rect 47961 11509 47995 11543
rect 47995 11509 48004 11543
rect 47952 11500 48004 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 47952 11228 48004 11280
rect 46664 11203 46716 11212
rect 46664 11169 46673 11203
rect 46673 11169 46707 11203
rect 46707 11169 46716 11203
rect 46664 11160 46716 11169
rect 46848 11160 46900 11212
rect 2964 11092 3016 11144
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2136 10004 2188 10056
rect 3148 10004 3200 10056
rect 41420 10004 41472 10056
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2872 9596 2924 9648
rect 41420 9596 41472 9648
rect 45192 9596 45244 9648
rect 47768 9596 47820 9648
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 2504 8916 2556 8968
rect 4620 8916 4672 8968
rect 2320 8780 2372 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2320 8551 2372 8560
rect 2320 8517 2329 8551
rect 2329 8517 2363 8551
rect 2363 8517 2372 8551
rect 2320 8508 2372 8517
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 44364 8440 44416 8492
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 41420 8415 41472 8424
rect 2780 8372 2832 8381
rect 41420 8381 41429 8415
rect 41429 8381 41463 8415
rect 41463 8381 41472 8415
rect 41420 8372 41472 8381
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 47492 7939 47544 7948
rect 47492 7905 47501 7939
rect 47501 7905 47535 7939
rect 47535 7905 47544 7939
rect 47492 7896 47544 7905
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 2412 7760 2464 7812
rect 5816 7828 5868 7880
rect 46020 7828 46072 7880
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4068 7420 4120 7472
rect 4620 7352 4672 7404
rect 24584 7352 24636 7404
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 5080 7327 5132 7336
rect 2780 7284 2832 7293
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 2964 7216 3016 7268
rect 1676 7148 1728 7200
rect 5080 7148 5132 7200
rect 47952 7191 48004 7200
rect 47952 7157 47961 7191
rect 47961 7157 47995 7191
rect 47995 7157 48004 7191
rect 47952 7148 48004 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6944 1636 6996
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 47952 6876 48004 6928
rect 48228 6851 48280 6860
rect 48228 6817 48237 6851
rect 48237 6817 48271 6851
rect 48271 6817 48280 6851
rect 48228 6808 48280 6817
rect 3056 6740 3108 6792
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 47860 6672 47912 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 47860 6443 47912 6452
rect 47860 6409 47869 6443
rect 47869 6409 47903 6443
rect 47903 6409 47912 6443
rect 47860 6400 47912 6409
rect 47584 6332 47636 6384
rect 47216 6264 47268 6316
rect 47400 6264 47452 6316
rect 48044 6264 48096 6316
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 2872 6196 2924 6248
rect 2964 6239 3016 6248
rect 2964 6205 2973 6239
rect 2973 6205 3007 6239
rect 3007 6205 3016 6239
rect 2964 6196 3016 6205
rect 4988 6060 5040 6112
rect 46480 6103 46532 6112
rect 46480 6069 46489 6103
rect 46489 6069 46523 6103
rect 46523 6069 46532 6103
rect 46480 6060 46532 6069
rect 46664 6060 46716 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2136 5856 2188 5908
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 3976 5788 4028 5840
rect 4712 5720 4764 5772
rect 17408 5720 17460 5772
rect 46664 5763 46716 5772
rect 46664 5729 46673 5763
rect 46673 5729 46707 5763
rect 46707 5729 46716 5763
rect 46664 5720 46716 5729
rect 48228 5763 48280 5772
rect 48228 5729 48237 5763
rect 48237 5729 48271 5763
rect 48271 5729 48280 5763
rect 48228 5720 48280 5729
rect 3792 5652 3844 5704
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 46020 5695 46072 5704
rect 46020 5661 46029 5695
rect 46029 5661 46063 5695
rect 46063 5661 46072 5695
rect 46020 5652 46072 5661
rect 10416 5584 10468 5636
rect 47952 5584 48004 5636
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4804 5312 4856 5364
rect 4068 5244 4120 5296
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 5724 5176 5776 5228
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 46020 5244 46072 5296
rect 5816 5176 5868 5185
rect 47952 5219 48004 5228
rect 47952 5185 47961 5219
rect 47961 5185 47995 5219
rect 47995 5185 48004 5219
rect 47952 5176 48004 5185
rect 2780 5108 2832 5117
rect 5080 5108 5132 5160
rect 8300 5108 8352 5160
rect 44548 5108 44600 5160
rect 48964 5108 49016 5160
rect 4804 4972 4856 5024
rect 4896 4972 4948 5024
rect 5632 4972 5684 5024
rect 44180 4972 44232 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 44548 4811 44600 4820
rect 44548 4777 44557 4811
rect 44557 4777 44591 4811
rect 44591 4777 44600 4811
rect 44548 4768 44600 4777
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 7012 4564 7064 4616
rect 40040 4564 40092 4616
rect 44272 4564 44324 4616
rect 48136 4700 48188 4752
rect 47952 4632 48004 4684
rect 45192 4607 45244 4616
rect 45192 4573 45201 4607
rect 45201 4573 45235 4607
rect 45235 4573 45244 4607
rect 45192 4564 45244 4573
rect 45744 4564 45796 4616
rect 1768 4539 1820 4548
rect 1768 4505 1777 4539
rect 1777 4505 1811 4539
rect 1811 4505 1820 4539
rect 1768 4496 1820 4505
rect 46480 4496 46532 4548
rect 48320 4539 48372 4548
rect 48320 4505 48329 4539
rect 48329 4505 48363 4539
rect 48363 4505 48372 4539
rect 48320 4496 48372 4505
rect 45376 4428 45428 4480
rect 45836 4428 45888 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 1768 4224 1820 4276
rect 1584 4088 1636 4140
rect 3148 4131 3200 4140
rect 1952 4020 2004 4072
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 8300 4131 8352 4140
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 10416 4131 10468 4140
rect 8300 4088 8352 4097
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 4068 3952 4120 4004
rect 10600 4020 10652 4072
rect 12900 4088 12952 4140
rect 20720 4020 20772 4072
rect 12900 3952 12952 4004
rect 44364 4131 44416 4140
rect 38660 4063 38712 4072
rect 38660 4029 38669 4063
rect 38669 4029 38703 4063
rect 38703 4029 38712 4063
rect 38660 4020 38712 4029
rect 39396 4020 39448 4072
rect 39304 3952 39356 4004
rect 44364 4097 44373 4131
rect 44373 4097 44407 4131
rect 44407 4097 44416 4131
rect 44364 4088 44416 4097
rect 47952 4131 48004 4140
rect 47952 4097 47961 4131
rect 47961 4097 47995 4131
rect 47995 4097 48004 4131
rect 47952 4088 48004 4097
rect 46940 4020 46992 4072
rect 47676 4020 47728 4072
rect 3976 3884 4028 3936
rect 6920 3884 6972 3936
rect 7564 3884 7616 3936
rect 8392 3927 8444 3936
rect 8392 3893 8401 3927
rect 8401 3893 8435 3927
rect 8435 3893 8444 3927
rect 8392 3884 8444 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 12532 3884 12584 3936
rect 13176 3884 13228 3936
rect 24768 3884 24820 3936
rect 25872 3884 25924 3936
rect 40500 3884 40552 3936
rect 42616 3884 42668 3936
rect 42984 3884 43036 3936
rect 45100 3884 45152 3936
rect 47952 3952 48004 4004
rect 47768 3884 47820 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4712 3680 4764 3732
rect 4804 3680 4856 3732
rect 5540 3680 5592 3732
rect 5356 3612 5408 3664
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 3148 3544 3200 3596
rect 3976 3544 4028 3596
rect 24584 3680 24636 3732
rect 44364 3680 44416 3732
rect 6460 3544 6512 3596
rect 10508 3587 10560 3596
rect 10508 3553 10517 3587
rect 10517 3553 10551 3587
rect 10551 3553 10560 3587
rect 10508 3544 10560 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 4160 3476 4212 3528
rect 10324 3519 10376 3528
rect 2596 3408 2648 3460
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 12992 3476 13044 3528
rect 16856 3476 16908 3528
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 19340 3476 19392 3528
rect 47032 3612 47084 3664
rect 25872 3587 25924 3596
rect 20260 3519 20312 3528
rect 20260 3485 20269 3519
rect 20269 3485 20303 3519
rect 20303 3485 20312 3519
rect 20260 3476 20312 3485
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 20720 3476 20772 3485
rect 22008 3476 22060 3528
rect 25872 3553 25881 3587
rect 25881 3553 25915 3587
rect 25915 3553 25924 3587
rect 25872 3544 25924 3553
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 39396 3587 39448 3596
rect 39396 3553 39405 3587
rect 39405 3553 39439 3587
rect 39439 3553 39448 3587
rect 39396 3544 39448 3553
rect 40500 3587 40552 3596
rect 40500 3553 40509 3587
rect 40509 3553 40543 3587
rect 40543 3553 40552 3587
rect 40500 3544 40552 3553
rect 41236 3587 41288 3596
rect 41236 3553 41245 3587
rect 41245 3553 41279 3587
rect 41279 3553 41288 3587
rect 41236 3544 41288 3553
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 27436 3476 27488 3528
rect 31852 3519 31904 3528
rect 31852 3485 31861 3519
rect 31861 3485 31895 3519
rect 31895 3485 31904 3519
rect 31852 3476 31904 3485
rect 32312 3519 32364 3528
rect 32312 3485 32321 3519
rect 32321 3485 32355 3519
rect 32355 3485 32364 3519
rect 32312 3476 32364 3485
rect 38384 3476 38436 3528
rect 17040 3340 17092 3392
rect 19432 3340 19484 3392
rect 20812 3383 20864 3392
rect 20812 3349 20821 3383
rect 20821 3349 20855 3383
rect 20855 3349 20864 3383
rect 20812 3340 20864 3349
rect 22192 3340 22244 3392
rect 24952 3340 25004 3392
rect 27528 3340 27580 3392
rect 32496 3340 32548 3392
rect 38568 3340 38620 3392
rect 42432 3476 42484 3528
rect 44272 3544 44324 3596
rect 44456 3476 44508 3528
rect 44916 3476 44968 3528
rect 41420 3408 41472 3460
rect 45836 3451 45888 3460
rect 42800 3340 42852 3392
rect 45836 3417 45845 3451
rect 45845 3417 45879 3451
rect 45879 3417 45888 3451
rect 45836 3408 45888 3417
rect 47032 3408 47084 3460
rect 47400 3340 47452 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4988 3136 5040 3188
rect 5632 3068 5684 3120
rect 8392 3068 8444 3120
rect 13176 3111 13228 3120
rect 13176 3077 13185 3111
rect 13185 3077 13219 3111
rect 13219 3077 13228 3111
rect 13176 3068 13228 3077
rect 17040 3111 17092 3120
rect 17040 3077 17049 3111
rect 17049 3077 17083 3111
rect 17083 3077 17092 3111
rect 17040 3068 17092 3077
rect 20812 3068 20864 3120
rect 22192 3111 22244 3120
rect 22192 3077 22201 3111
rect 22201 3077 22235 3111
rect 22235 3077 22244 3111
rect 22192 3068 22244 3077
rect 24952 3111 25004 3120
rect 24952 3077 24961 3111
rect 24961 3077 24995 3111
rect 24995 3077 25004 3111
rect 24952 3068 25004 3077
rect 32496 3111 32548 3120
rect 32496 3077 32505 3111
rect 32505 3077 32539 3111
rect 32539 3077 32548 3111
rect 32496 3068 32548 3077
rect 38568 3111 38620 3120
rect 38568 3077 38577 3111
rect 38577 3077 38611 3111
rect 38611 3077 38620 3111
rect 38568 3068 38620 3077
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 10324 3000 10376 3052
rect 10600 3000 10652 3052
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 31852 3000 31904 3052
rect 38384 3043 38436 3052
rect 38384 3009 38393 3043
rect 38393 3009 38427 3043
rect 38427 3009 38436 3043
rect 38384 3000 38436 3009
rect 45744 3136 45796 3188
rect 41420 3111 41472 3120
rect 41420 3077 41429 3111
rect 41429 3077 41463 3111
rect 41463 3077 41472 3111
rect 41420 3068 41472 3077
rect 42800 3111 42852 3120
rect 42800 3077 42809 3111
rect 42809 3077 42843 3111
rect 42843 3077 42852 3111
rect 42800 3068 42852 3077
rect 45100 3111 45152 3120
rect 45100 3077 45109 3111
rect 45109 3077 45143 3111
rect 45143 3077 45152 3111
rect 45100 3068 45152 3077
rect 42432 3000 42484 3052
rect 42616 3043 42668 3052
rect 42616 3009 42625 3043
rect 42625 3009 42659 3043
rect 42659 3009 42668 3043
rect 42616 3000 42668 3009
rect 44916 3043 44968 3052
rect 44916 3009 44925 3043
rect 44925 3009 44959 3043
rect 44959 3009 44968 3043
rect 44916 3000 44968 3009
rect 47952 3043 48004 3052
rect 47952 3009 47961 3043
rect 47961 3009 47995 3043
rect 47995 3009 48004 3043
rect 47952 3000 48004 3009
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7840 2932 7892 2984
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 20260 2932 20312 2984
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 25780 2975 25832 2984
rect 25780 2941 25789 2975
rect 25789 2941 25823 2975
rect 25823 2941 25832 2975
rect 25780 2932 25832 2941
rect 27620 2975 27672 2984
rect 27620 2941 27629 2975
rect 27629 2941 27663 2975
rect 27663 2941 27672 2975
rect 27620 2932 27672 2941
rect 27712 2932 27764 2984
rect 32220 2932 32272 2984
rect 4712 2864 4764 2916
rect 41880 2932 41932 2984
rect 45100 2932 45152 2984
rect 46756 2864 46808 2916
rect 3240 2796 3292 2848
rect 4068 2796 4120 2848
rect 7104 2839 7156 2848
rect 7104 2805 7113 2839
rect 7113 2805 7147 2839
rect 7147 2805 7156 2839
rect 7104 2796 7156 2805
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 40224 2796 40276 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3792 2592 3844 2644
rect 4712 2635 4764 2644
rect 4712 2601 4721 2635
rect 4721 2601 4755 2635
rect 4755 2601 4764 2635
rect 5632 2635 5684 2644
rect 4712 2592 4764 2601
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 5724 2524 5776 2576
rect 12900 2592 12952 2644
rect 27620 2635 27672 2644
rect 27620 2601 27629 2635
rect 27629 2601 27663 2635
rect 27663 2601 27672 2635
rect 27620 2592 27672 2601
rect 38660 2592 38712 2644
rect 46940 2592 46992 2644
rect 664 2456 716 2508
rect 7104 2456 7156 2508
rect 7196 2499 7248 2508
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 12532 2524 12584 2576
rect 19432 2524 19484 2576
rect 7196 2456 7248 2465
rect 12440 2456 12492 2508
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 19708 2456 19760 2508
rect 24308 2456 24360 2508
rect 40040 2499 40092 2508
rect 40040 2465 40049 2499
rect 40049 2465 40083 2499
rect 40083 2465 40092 2499
rect 40040 2456 40092 2465
rect 40224 2499 40276 2508
rect 40224 2465 40233 2499
rect 40233 2465 40267 2499
rect 40267 2465 40276 2499
rect 40224 2456 40276 2465
rect 40592 2499 40644 2508
rect 40592 2465 40601 2499
rect 40601 2465 40635 2499
rect 40635 2465 40644 2499
rect 40592 2456 40644 2465
rect 44180 2524 44232 2576
rect 42984 2499 43036 2508
rect 42984 2465 42993 2499
rect 42993 2465 43027 2499
rect 43027 2465 43036 2499
rect 42984 2456 43036 2465
rect 44456 2456 44508 2508
rect 45376 2499 45428 2508
rect 45376 2465 45385 2499
rect 45385 2465 45419 2499
rect 45419 2465 45428 2499
rect 45376 2456 45428 2465
rect 45744 2499 45796 2508
rect 45744 2465 45753 2499
rect 45753 2465 45787 2499
rect 45787 2465 45796 2499
rect 45744 2456 45796 2465
rect 4160 2388 4212 2440
rect 5724 2388 5776 2440
rect 19340 2388 19392 2440
rect 23848 2388 23900 2440
rect 27528 2431 27580 2440
rect 27528 2397 27537 2431
rect 27537 2397 27571 2431
rect 27571 2397 27580 2431
rect 27528 2388 27580 2397
rect 32312 2388 32364 2440
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 4896 2320 4948 2372
rect 6920 2363 6972 2372
rect 6920 2329 6929 2363
rect 6929 2329 6963 2363
rect 6963 2329 6972 2363
rect 6920 2320 6972 2329
rect 7012 2252 7064 2304
rect 46848 2252 46900 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect -10 49200 102 49800
rect 1278 49200 1390 49800
rect 1922 49200 2034 49800
rect 2566 49200 2678 49800
rect 3854 49200 3966 49800
rect 4498 49314 4610 49800
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 32 48822 60 49200
rect 20 48816 72 48822
rect 20 48758 72 48764
rect 1768 46912 1820 46918
rect 1768 46854 1820 46860
rect 1780 46034 1808 46854
rect 1964 46442 1992 49200
rect 2044 47048 2096 47054
rect 2044 46990 2096 46996
rect 1952 46436 2004 46442
rect 1952 46378 2004 46384
rect 1768 46028 1820 46034
rect 1768 45970 1820 45976
rect 2056 45554 2084 46990
rect 2608 46510 2636 49200
rect 2778 48376 2834 48385
rect 2778 48311 2834 48320
rect 2688 47048 2740 47054
rect 2688 46990 2740 46996
rect 2596 46504 2648 46510
rect 2596 46446 2648 46452
rect 1964 45526 2084 45554
rect 1768 44872 1820 44878
rect 1768 44814 1820 44820
rect 1584 43784 1636 43790
rect 1584 43726 1636 43732
rect 1596 43314 1624 43726
rect 1584 43308 1636 43314
rect 1584 43250 1636 43256
rect 1780 26234 1808 44814
rect 1964 43246 1992 45526
rect 2504 45416 2556 45422
rect 2504 45358 2556 45364
rect 2320 45348 2372 45354
rect 2320 45290 2372 45296
rect 2228 45280 2280 45286
rect 2228 45222 2280 45228
rect 2240 44402 2268 45222
rect 2228 44396 2280 44402
rect 2228 44338 2280 44344
rect 1952 43240 2004 43246
rect 1952 43182 2004 43188
rect 1688 26206 1808 26234
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25362 1624 25638
rect 1584 25356 1636 25362
rect 1584 25298 1636 25304
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21554 1624 21966
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13938 1624 14350
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7002 1624 7822
rect 1688 7206 1716 26206
rect 1768 25220 1820 25226
rect 1768 25162 1820 25168
rect 1780 24954 1808 25162
rect 1768 24948 1820 24954
rect 1768 24890 1820 24896
rect 1768 21956 1820 21962
rect 1768 21898 1820 21904
rect 1780 21690 1808 21898
rect 1768 21684 1820 21690
rect 1768 21626 1820 21632
rect 1964 16574 1992 43182
rect 2332 42770 2360 45290
rect 2412 44736 2464 44742
rect 2412 44678 2464 44684
rect 2424 44470 2452 44678
rect 2516 44538 2544 45358
rect 2504 44532 2556 44538
rect 2504 44474 2556 44480
rect 2412 44464 2464 44470
rect 2412 44406 2464 44412
rect 2596 43716 2648 43722
rect 2596 43658 2648 43664
rect 2608 43450 2636 43658
rect 2596 43444 2648 43450
rect 2596 43386 2648 43392
rect 2320 42764 2372 42770
rect 2320 42706 2372 42712
rect 2700 42566 2728 46990
rect 2792 46034 2820 48311
rect 3514 47696 3570 47705
rect 3514 47631 3570 47640
rect 3528 47122 3556 47631
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 3516 47116 3568 47122
rect 3516 47058 3568 47064
rect 4160 47048 4212 47054
rect 4160 46990 4212 46996
rect 4068 46640 4120 46646
rect 4068 46582 4120 46588
rect 2964 46436 3016 46442
rect 2964 46378 3016 46384
rect 2870 46336 2926 46345
rect 2870 46271 2926 46280
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2778 45656 2834 45665
rect 2778 45591 2834 45600
rect 2792 44334 2820 45591
rect 2780 44328 2832 44334
rect 2780 44270 2832 44276
rect 2780 43852 2832 43858
rect 2780 43794 2832 43800
rect 2792 43625 2820 43794
rect 2778 43616 2834 43625
rect 2778 43551 2834 43560
rect 2884 42702 2912 46271
rect 2976 45422 3004 46378
rect 3056 45892 3108 45898
rect 3056 45834 3108 45840
rect 2964 45416 3016 45422
rect 2964 45358 3016 45364
rect 3068 42770 3096 45834
rect 3240 44804 3292 44810
rect 3240 44746 3292 44752
rect 3056 42764 3108 42770
rect 3056 42706 3108 42712
rect 2872 42696 2924 42702
rect 2872 42638 2924 42644
rect 2688 42560 2740 42566
rect 2688 42502 2740 42508
rect 2044 41608 2096 41614
rect 2044 41550 2096 41556
rect 2056 41138 2084 41550
rect 2044 41132 2096 41138
rect 2044 41074 2096 41080
rect 2412 41064 2464 41070
rect 2412 41006 2464 41012
rect 2780 41064 2832 41070
rect 2780 41006 2832 41012
rect 2424 40730 2452 41006
rect 2792 40905 2820 41006
rect 2778 40896 2834 40905
rect 2778 40831 2834 40840
rect 2412 40724 2464 40730
rect 2412 40666 2464 40672
rect 2228 40520 2280 40526
rect 2228 40462 2280 40468
rect 2240 26234 2268 40462
rect 2320 33312 2372 33318
rect 2320 33254 2372 33260
rect 2332 32978 2360 33254
rect 2320 32972 2372 32978
rect 2320 32914 2372 32920
rect 2780 32972 2832 32978
rect 2780 32914 2832 32920
rect 2412 32836 2464 32842
rect 2412 32778 2464 32784
rect 2424 32570 2452 32778
rect 2792 32745 2820 32914
rect 2778 32736 2834 32745
rect 2778 32671 2834 32680
rect 2412 32564 2464 32570
rect 2412 32506 2464 32512
rect 2596 32428 2648 32434
rect 2596 32370 2648 32376
rect 2240 26206 2360 26234
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 2056 23730 2084 24142
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 2240 23322 2268 23598
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 2332 21418 2360 26206
rect 2412 23112 2464 23118
rect 2412 23054 2464 23060
rect 2424 22710 2452 23054
rect 2412 22704 2464 22710
rect 2412 22646 2464 22652
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 2056 20466 2084 20878
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2056 18290 2084 18702
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2056 16794 2084 17070
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 1964 16546 2084 16574
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1964 15026 1992 15438
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1780 14074 1808 14282
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 2056 6914 2084 16546
rect 2148 15502 2176 19790
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2240 17882 2268 18158
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2240 15094 2268 15302
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2332 11830 2360 12174
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2332 11354 2360 11630
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9586 2176 9998
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8498 2176 8910
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8566 2360 8774
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2424 7818 2452 22646
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2516 20058 2544 20334
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2516 8974 2544 17614
rect 2608 16658 2636 32370
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2792 25265 2820 25298
rect 2778 25256 2834 25265
rect 2778 25191 2834 25200
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2778 23896 2834 23905
rect 2778 23831 2834 23840
rect 2792 23662 2820 23831
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 2792 21865 2820 22034
rect 2778 21856 2834 21865
rect 2778 21791 2834 21800
rect 2976 21554 3004 24754
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 2688 21412 2740 21418
rect 2688 21354 2740 21360
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 1964 6886 2084 6914
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 4146 1624 4558
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1780 4282 1808 4490
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1964 4078 1992 6886
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2148 5914 2176 6190
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 2608 3466 2636 15438
rect 2700 13938 2728 21354
rect 2778 20496 2834 20505
rect 2778 20431 2834 20440
rect 2792 20398 2820 20431
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 18222 2820 18391
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2780 17128 2832 17134
rect 2778 17096 2780 17105
rect 2832 17096 2834 17105
rect 2778 17031 2834 17040
rect 2884 16522 2912 17206
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14385 2820 14418
rect 2778 14376 2834 14385
rect 2778 14311 2834 14320
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2976 11150 3004 21490
rect 3252 19854 3280 44746
rect 3976 44260 4028 44266
rect 3976 44202 4028 44208
rect 3988 43790 4016 44202
rect 4080 43994 4108 46582
rect 4172 46578 4200 46990
rect 4160 46572 4212 46578
rect 4160 46514 4212 46520
rect 4724 46510 4752 49286
rect 5786 49200 5898 49800
rect 6430 49200 6542 49800
rect 7718 49200 7830 49800
rect 8362 49200 8474 49800
rect 9006 49200 9118 49800
rect 10294 49200 10406 49800
rect 10938 49200 11050 49800
rect 12226 49200 12338 49800
rect 12870 49200 12982 49800
rect 14158 49200 14270 49800
rect 14802 49200 14914 49800
rect 15446 49200 15558 49800
rect 16734 49200 16846 49800
rect 17378 49200 17490 49800
rect 18666 49200 18778 49800
rect 19310 49200 19422 49800
rect 20598 49200 20710 49800
rect 21242 49200 21354 49800
rect 21886 49200 21998 49800
rect 23174 49200 23286 49800
rect 23818 49200 23930 49800
rect 25106 49200 25218 49800
rect 25750 49200 25862 49800
rect 27038 49200 27150 49800
rect 27682 49314 27794 49800
rect 27682 49286 28028 49314
rect 27682 49200 27794 49286
rect 4896 47184 4948 47190
rect 4896 47126 4948 47132
rect 4804 46980 4856 46986
rect 4804 46922 4856 46928
rect 4620 46504 4672 46510
rect 4620 46446 4672 46452
rect 4712 46504 4764 46510
rect 4712 46446 4764 46452
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4632 45082 4660 46446
rect 4816 45966 4844 46922
rect 4908 46170 4936 47126
rect 5540 47048 5592 47054
rect 5540 46990 5592 46996
rect 5724 47048 5776 47054
rect 5724 46990 5776 46996
rect 4896 46164 4948 46170
rect 4896 46106 4948 46112
rect 4908 46034 4936 46106
rect 5552 46034 5580 46990
rect 4896 46028 4948 46034
rect 4896 45970 4948 45976
rect 5540 46028 5592 46034
rect 5540 45970 5592 45976
rect 4804 45960 4856 45966
rect 4804 45902 4856 45908
rect 4816 45554 4844 45902
rect 4724 45526 4844 45554
rect 4724 45490 4752 45526
rect 4712 45484 4764 45490
rect 4712 45426 4764 45432
rect 4896 45484 4948 45490
rect 4896 45426 4948 45432
rect 4620 45076 4672 45082
rect 4620 45018 4672 45024
rect 4724 44742 4752 45426
rect 4908 44878 4936 45426
rect 4988 45416 5040 45422
rect 4988 45358 5040 45364
rect 4896 44872 4948 44878
rect 4896 44814 4948 44820
rect 4528 44736 4580 44742
rect 4528 44678 4580 44684
rect 4712 44736 4764 44742
rect 4712 44678 4764 44684
rect 4540 44402 4568 44678
rect 4528 44396 4580 44402
rect 4528 44338 4580 44344
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4068 43988 4120 43994
rect 4068 43930 4120 43936
rect 4724 43790 4752 44678
rect 5000 43858 5028 45358
rect 5736 44810 5764 46990
rect 5828 46034 5856 49200
rect 8024 48816 8076 48822
rect 8024 48758 8076 48764
rect 7012 47116 7064 47122
rect 7012 47058 7064 47064
rect 6552 47048 6604 47054
rect 6552 46990 6604 46996
rect 6564 46578 6592 46990
rect 6736 46912 6788 46918
rect 6736 46854 6788 46860
rect 6748 46646 6776 46854
rect 6736 46640 6788 46646
rect 6736 46582 6788 46588
rect 6552 46572 6604 46578
rect 6552 46514 6604 46520
rect 7024 46510 7052 47058
rect 8036 47054 8064 48758
rect 8404 47054 8432 49200
rect 7380 47048 7432 47054
rect 7380 46990 7432 46996
rect 8024 47048 8076 47054
rect 8024 46990 8076 46996
rect 8392 47048 8444 47054
rect 8392 46990 8444 46996
rect 7392 46714 7420 46990
rect 7840 46912 7892 46918
rect 7840 46854 7892 46860
rect 9128 46912 9180 46918
rect 9128 46854 9180 46860
rect 7380 46708 7432 46714
rect 7380 46650 7432 46656
rect 7012 46504 7064 46510
rect 7012 46446 7064 46452
rect 5816 46028 5868 46034
rect 5816 45970 5868 45976
rect 6644 45892 6696 45898
rect 6644 45834 6696 45840
rect 6656 45626 6684 45834
rect 6644 45620 6696 45626
rect 6644 45562 6696 45568
rect 5724 44804 5776 44810
rect 5724 44746 5776 44752
rect 5448 44328 5500 44334
rect 5448 44270 5500 44276
rect 4988 43852 5040 43858
rect 4988 43794 5040 43800
rect 3976 43784 4028 43790
rect 3976 43726 4028 43732
rect 4712 43784 4764 43790
rect 4712 43726 4764 43732
rect 3514 41576 3570 41585
rect 3514 41511 3570 41520
rect 3528 23798 3556 41511
rect 3988 24818 4016 43726
rect 4620 43444 4672 43450
rect 4620 43386 4672 43392
rect 4632 43246 4660 43386
rect 4724 43314 4752 43726
rect 4712 43308 4764 43314
rect 4712 43250 4764 43256
rect 4620 43240 4672 43246
rect 4620 43182 4672 43188
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3516 23792 3568 23798
rect 3516 23734 3568 23740
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17678 4660 43182
rect 4724 42922 4752 43250
rect 4724 42894 4844 42922
rect 4712 42764 4764 42770
rect 4712 42706 4764 42712
rect 4724 42294 4752 42706
rect 4816 42702 4844 42894
rect 4804 42696 4856 42702
rect 4804 42638 4856 42644
rect 4712 42288 4764 42294
rect 4712 42230 4764 42236
rect 4724 40526 4752 42230
rect 4712 40520 4764 40526
rect 4712 40462 4764 40468
rect 5460 22710 5488 44270
rect 5540 43852 5592 43858
rect 5540 43794 5592 43800
rect 5552 43722 5580 43794
rect 5540 43716 5592 43722
rect 5540 43658 5592 43664
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2962 10296 3018 10305
rect 2962 10231 3018 10240
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9654 2912 9862
rect 2872 9648 2924 9654
rect 2778 9616 2834 9625
rect 2872 9590 2924 9596
rect 2778 9551 2834 9560
rect 2792 8430 2820 9551
rect 2976 9518 3004 10231
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7585 3004 7890
rect 2962 7576 3018 7585
rect 2962 7511 3018 7520
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2792 6905 2820 7278
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2778 6896 2834 6905
rect 2976 6866 3004 7210
rect 2778 6831 2834 6840
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3068 6798 3096 13874
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2884 5914 2912 6190
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2976 5545 3004 6190
rect 2962 5536 3018 5545
rect 2962 5471 3018 5480
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4865 2820 5102
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2792 2825 2820 3538
rect 2976 3505 3004 4626
rect 3160 4146 3188 9998
rect 3804 5710 3832 16594
rect 5552 16574 5580 43658
rect 5552 16546 5672 16574
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4080 6866 4108 7414
rect 4632 7410 4660 8910
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5092 7206 5120 7278
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 5846 4016 6734
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5302 4108 5510
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3160 3602 3188 4082
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 2962 3496 3018 3505
rect 2962 3431 3018 3440
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 664 2508 716 2514
rect 664 2450 716 2456
rect 676 800 704 2450
rect 2884 1465 2912 2926
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3252 800 3280 2790
rect 3804 2650 3832 4014
rect 3988 3942 4016 4014
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3988 2666 4016 3538
rect 4080 2854 4108 3946
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4724 3738 4752 5714
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 5370 4844 5646
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4816 3890 4844 4966
rect 4908 4690 4936 4966
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4816 3862 4936 3890
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 3058 4200 3470
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3792 2644 3844 2650
rect 3988 2638 4108 2666
rect 4724 2650 4752 2858
rect 3792 2586 3844 2592
rect 4080 2530 4108 2638
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4080 2502 4200 2530
rect 4172 2446 4200 2502
rect 4160 2440 4212 2446
rect 4816 2394 4844 3674
rect 4160 2382 4212 2388
rect 4540 2366 4844 2394
rect 4908 2378 4936 3862
rect 5000 3194 5028 6054
rect 5092 5166 5120 7142
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5644 5114 5672 16546
rect 5736 5234 5764 44746
rect 7380 44464 7432 44470
rect 7380 44406 7432 44412
rect 7392 32434 7420 44406
rect 7852 43382 7880 46854
rect 7840 43376 7892 43382
rect 7840 43318 7892 43324
rect 9140 43314 9168 46854
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 46034 10456 46310
rect 10980 46034 11008 49200
rect 12532 47048 12584 47054
rect 12532 46990 12584 46996
rect 12544 46646 12572 46990
rect 12532 46640 12584 46646
rect 12532 46582 12584 46588
rect 12912 46510 12940 49200
rect 12440 46504 12492 46510
rect 12440 46446 12492 46452
rect 12900 46504 12952 46510
rect 12900 46446 12952 46452
rect 10416 46028 10468 46034
rect 10416 45970 10468 45976
rect 10968 46028 11020 46034
rect 10968 45970 11020 45976
rect 10600 45892 10652 45898
rect 10600 45834 10652 45840
rect 10612 45626 10640 45834
rect 10600 45620 10652 45626
rect 10600 45562 10652 45568
rect 12452 45558 12480 46446
rect 13360 45960 13412 45966
rect 13360 45902 13412 45908
rect 13544 45960 13596 45966
rect 13544 45902 13596 45908
rect 12440 45552 12492 45558
rect 12440 45494 12492 45500
rect 13372 45490 13400 45902
rect 13556 45626 13584 45902
rect 13544 45620 13596 45626
rect 13544 45562 13596 45568
rect 10508 45484 10560 45490
rect 10508 45426 10560 45432
rect 12348 45484 12400 45490
rect 12348 45426 12400 45432
rect 12992 45484 13044 45490
rect 12992 45426 13044 45432
rect 13360 45484 13412 45490
rect 13360 45426 13412 45432
rect 10324 45416 10376 45422
rect 10520 45370 10548 45426
rect 10376 45364 10548 45370
rect 10324 45358 10548 45364
rect 10336 45342 10548 45358
rect 9128 43308 9180 43314
rect 9128 43250 9180 43256
rect 10520 32502 10548 45342
rect 12360 45286 12388 45426
rect 12348 45280 12400 45286
rect 12348 45222 12400 45228
rect 12360 44810 12388 45222
rect 12348 44804 12400 44810
rect 12348 44746 12400 44752
rect 13004 44470 13032 45426
rect 12992 44464 13044 44470
rect 12992 44406 13044 44412
rect 10508 32496 10560 32502
rect 10508 32438 10560 32444
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 13004 28218 13032 44406
rect 13556 43722 13584 45562
rect 14200 45422 14228 49200
rect 14556 47048 14608 47054
rect 14556 46990 14608 46996
rect 14568 46034 14596 46990
rect 14648 46504 14700 46510
rect 14648 46446 14700 46452
rect 14660 46102 14688 46446
rect 14648 46096 14700 46102
rect 14648 46038 14700 46044
rect 14844 46034 14872 49200
rect 15200 47048 15252 47054
rect 15200 46990 15252 46996
rect 15212 46646 15240 46990
rect 15200 46640 15252 46646
rect 15200 46582 15252 46588
rect 15488 46510 15516 49200
rect 22468 47048 22520 47054
rect 22468 46990 22520 46996
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 22480 46578 22508 46990
rect 22468 46572 22520 46578
rect 22468 46514 22520 46520
rect 23216 46510 23244 49200
rect 15476 46504 15528 46510
rect 15476 46446 15528 46452
rect 22928 46504 22980 46510
rect 22928 46446 22980 46452
rect 23204 46504 23256 46510
rect 23204 46446 23256 46452
rect 24952 46504 25004 46510
rect 24952 46446 25004 46452
rect 22744 46368 22796 46374
rect 22744 46310 22796 46316
rect 22756 46170 22784 46310
rect 22940 46170 22968 46446
rect 22744 46164 22796 46170
rect 22744 46106 22796 46112
rect 22928 46164 22980 46170
rect 22928 46106 22980 46112
rect 14556 46028 14608 46034
rect 14556 45970 14608 45976
rect 14832 46028 14884 46034
rect 14832 45970 14884 45976
rect 16580 45960 16632 45966
rect 16580 45902 16632 45908
rect 14188 45416 14240 45422
rect 14188 45358 14240 45364
rect 16592 45286 16620 45902
rect 24768 45892 24820 45898
rect 24768 45834 24820 45840
rect 22836 45824 22888 45830
rect 22836 45766 22888 45772
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 16580 45280 16632 45286
rect 16580 45222 16632 45228
rect 22848 44946 22876 45766
rect 24780 45626 24808 45834
rect 24964 45626 24992 46446
rect 25148 46034 25176 49200
rect 25320 47048 25372 47054
rect 25320 46990 25372 46996
rect 25332 46646 25360 46990
rect 25320 46640 25372 46646
rect 25320 46582 25372 46588
rect 25792 46510 25820 49200
rect 25780 46504 25832 46510
rect 25780 46446 25832 46452
rect 26976 46504 27028 46510
rect 26976 46446 27028 46452
rect 26988 46170 27016 46446
rect 27080 46442 27108 49200
rect 28000 47054 28028 49286
rect 28970 49200 29082 49800
rect 29614 49200 29726 49800
rect 30258 49200 30370 49800
rect 31546 49200 31658 49800
rect 32190 49200 32302 49800
rect 33478 49200 33590 49800
rect 34122 49200 34234 49800
rect 35410 49200 35522 49800
rect 36054 49200 36166 49800
rect 36698 49200 36810 49800
rect 37986 49200 38098 49800
rect 38630 49200 38742 49800
rect 39918 49200 40030 49800
rect 40562 49200 40674 49800
rect 41850 49200 41962 49800
rect 42494 49200 42606 49800
rect 43138 49200 43250 49800
rect 44426 49200 44538 49800
rect 45070 49200 45182 49800
rect 46358 49314 46470 49800
rect 45848 49286 46470 49314
rect 27160 47048 27212 47054
rect 27160 46990 27212 46996
rect 27988 47048 28040 47054
rect 27988 46990 28040 46996
rect 29092 47048 29144 47054
rect 29092 46990 29144 46996
rect 27172 46578 27200 46990
rect 27804 46912 27856 46918
rect 27804 46854 27856 46860
rect 27160 46572 27212 46578
rect 27160 46514 27212 46520
rect 27068 46436 27120 46442
rect 27068 46378 27120 46384
rect 26976 46164 27028 46170
rect 26976 46106 27028 46112
rect 25136 46028 25188 46034
rect 25136 45970 25188 45976
rect 26976 45960 27028 45966
rect 26976 45902 27028 45908
rect 24768 45620 24820 45626
rect 24768 45562 24820 45568
rect 24952 45620 25004 45626
rect 24952 45562 25004 45568
rect 26988 45354 27016 45902
rect 26976 45348 27028 45354
rect 26976 45290 27028 45296
rect 22836 44940 22888 44946
rect 22836 44882 22888 44888
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 13544 43716 13596 43722
rect 13544 43658 13596 43664
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 22376 43376 22428 43382
rect 22428 43324 22600 43330
rect 22376 43318 22600 43324
rect 22388 43314 22600 43318
rect 22388 43308 22612 43314
rect 22388 43302 22560 43308
rect 22560 43250 22612 43256
rect 23664 43172 23716 43178
rect 23664 43114 23716 43120
rect 23572 43104 23624 43110
rect 23572 43046 23624 43052
rect 23480 42560 23532 42566
rect 23480 42502 23532 42508
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 23492 42294 23520 42502
rect 23480 42288 23532 42294
rect 23480 42230 23532 42236
rect 23584 42226 23612 43046
rect 23676 42702 23704 43114
rect 23664 42696 23716 42702
rect 23664 42638 23716 42644
rect 23572 42220 23624 42226
rect 23572 42162 23624 42168
rect 24308 42220 24360 42226
rect 24308 42162 24360 42168
rect 23388 42016 23440 42022
rect 23388 41958 23440 41964
rect 23400 41546 23428 41958
rect 24320 41614 24348 42162
rect 24308 41608 24360 41614
rect 24308 41550 24360 41556
rect 23388 41540 23440 41546
rect 23388 41482 23440 41488
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 24320 41138 24348 41550
rect 24308 41132 24360 41138
rect 24308 41074 24360 41080
rect 24492 41132 24544 41138
rect 24492 41074 24544 41080
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 23940 40044 23992 40050
rect 23940 39986 23992 39992
rect 23952 39642 23980 39986
rect 24320 39846 24348 41074
rect 24504 40730 24532 41074
rect 25596 40928 25648 40934
rect 25596 40870 25648 40876
rect 24492 40724 24544 40730
rect 24492 40666 24544 40672
rect 24768 40520 24820 40526
rect 24768 40462 24820 40468
rect 24780 39982 24808 40462
rect 25044 40452 25096 40458
rect 25044 40394 25096 40400
rect 25056 40186 25084 40394
rect 25044 40180 25096 40186
rect 25044 40122 25096 40128
rect 24768 39976 24820 39982
rect 24768 39918 24820 39924
rect 24308 39840 24360 39846
rect 24308 39782 24360 39788
rect 24584 39840 24636 39846
rect 24584 39782 24636 39788
rect 23940 39636 23992 39642
rect 23940 39578 23992 39584
rect 24596 39574 24624 39782
rect 24584 39568 24636 39574
rect 24584 39510 24636 39516
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 23848 38208 23900 38214
rect 23848 38150 23900 38156
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 23860 37942 23888 38150
rect 23848 37936 23900 37942
rect 23848 37878 23900 37884
rect 24596 37874 24624 39510
rect 24780 39438 24808 39918
rect 24768 39432 24820 39438
rect 24688 39392 24768 39420
rect 24584 37868 24636 37874
rect 24584 37810 24636 37816
rect 23388 37120 23440 37126
rect 23388 37062 23440 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 23400 36174 23428 37062
rect 24032 36576 24084 36582
rect 24032 36518 24084 36524
rect 24044 36174 24072 36518
rect 23388 36168 23440 36174
rect 23388 36110 23440 36116
rect 24032 36168 24084 36174
rect 24032 36110 24084 36116
rect 23756 36032 23808 36038
rect 23756 35974 23808 35980
rect 24032 36032 24084 36038
rect 24032 35974 24084 35980
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 23768 35766 23796 35974
rect 23756 35760 23808 35766
rect 23756 35702 23808 35708
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 24044 34610 24072 35974
rect 24596 35630 24624 37810
rect 24688 37262 24716 39392
rect 24768 39374 24820 39380
rect 25056 39030 25084 40122
rect 25608 40050 25636 40870
rect 25596 40044 25648 40050
rect 25596 39986 25648 39992
rect 25608 39522 25636 39986
rect 26608 39840 26660 39846
rect 26608 39782 26660 39788
rect 25608 39494 25820 39522
rect 25596 39296 25648 39302
rect 25596 39238 25648 39244
rect 25688 39296 25740 39302
rect 25688 39238 25740 39244
rect 25608 39030 25636 39238
rect 25700 39098 25728 39238
rect 25792 39098 25820 39494
rect 26424 39364 26476 39370
rect 26424 39306 26476 39312
rect 26436 39098 26464 39306
rect 25688 39092 25740 39098
rect 25688 39034 25740 39040
rect 25780 39092 25832 39098
rect 25780 39034 25832 39040
rect 26424 39092 26476 39098
rect 26424 39034 26476 39040
rect 25044 39024 25096 39030
rect 25044 38966 25096 38972
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 25056 38350 25084 38966
rect 25608 38554 25636 38966
rect 25596 38548 25648 38554
rect 25596 38490 25648 38496
rect 24768 38344 24820 38350
rect 24768 38286 24820 38292
rect 25044 38344 25096 38350
rect 25044 38286 25096 38292
rect 24780 37466 24808 38286
rect 25608 38010 25636 38490
rect 25700 38418 25728 39034
rect 25688 38412 25740 38418
rect 25688 38354 25740 38360
rect 25792 38298 25820 39034
rect 26620 38962 26648 39782
rect 26608 38956 26660 38962
rect 26608 38898 26660 38904
rect 25964 38752 26016 38758
rect 25964 38694 26016 38700
rect 25700 38282 25820 38298
rect 25688 38276 25820 38282
rect 25740 38270 25820 38276
rect 25688 38218 25740 38224
rect 25596 38004 25648 38010
rect 25596 37946 25648 37952
rect 24768 37460 24820 37466
rect 24768 37402 24820 37408
rect 25320 37392 25372 37398
rect 25320 37334 25372 37340
rect 24952 37324 25004 37330
rect 24952 37266 25004 37272
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 24688 36786 24716 37198
rect 24964 36854 24992 37266
rect 24952 36848 25004 36854
rect 24952 36790 25004 36796
rect 24676 36780 24728 36786
rect 24676 36722 24728 36728
rect 25332 35698 25360 37334
rect 25976 36922 26004 38694
rect 26240 38208 26292 38214
rect 26240 38150 26292 38156
rect 26252 37398 26280 38150
rect 26056 37392 26108 37398
rect 26240 37392 26292 37398
rect 26108 37340 26188 37346
rect 26056 37334 26188 37340
rect 26240 37334 26292 37340
rect 26068 37318 26188 37334
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 25964 36916 26016 36922
rect 25964 36858 26016 36864
rect 25780 36848 25832 36854
rect 25780 36790 25832 36796
rect 25792 36666 25820 36790
rect 25792 36638 25912 36666
rect 26068 36650 26096 37198
rect 26160 36854 26188 37318
rect 26332 37256 26384 37262
rect 26332 37198 26384 37204
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 26252 36854 26280 37062
rect 26148 36848 26200 36854
rect 26148 36790 26200 36796
rect 26240 36848 26292 36854
rect 26240 36790 26292 36796
rect 25884 36582 25912 36638
rect 26056 36644 26108 36650
rect 26056 36586 26108 36592
rect 25780 36576 25832 36582
rect 25780 36518 25832 36524
rect 25872 36576 25924 36582
rect 26068 36530 26096 36586
rect 25872 36518 25924 36524
rect 25320 35692 25372 35698
rect 25320 35634 25372 35640
rect 24584 35624 24636 35630
rect 24584 35566 24636 35572
rect 24596 35086 24624 35566
rect 24584 35080 24636 35086
rect 24584 35022 24636 35028
rect 24596 34678 24624 35022
rect 25332 34746 25360 35634
rect 25792 35018 25820 36518
rect 25976 36502 26096 36530
rect 25976 35834 26004 36502
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26252 35850 26280 35974
rect 25964 35828 26016 35834
rect 25964 35770 26016 35776
rect 26068 35822 26280 35850
rect 25780 35012 25832 35018
rect 25780 34954 25832 34960
rect 26068 34950 26096 35822
rect 26344 35290 26372 37198
rect 26608 37188 26660 37194
rect 26608 37130 26660 37136
rect 26620 36718 26648 37130
rect 26988 36854 27016 45290
rect 27816 43790 27844 46854
rect 29104 46578 29132 46990
rect 29656 46594 29684 49200
rect 29920 47048 29972 47054
rect 29920 46990 29972 46996
rect 29092 46572 29144 46578
rect 29656 46566 29776 46594
rect 29092 46514 29144 46520
rect 29748 46510 29776 46566
rect 29644 46504 29696 46510
rect 29644 46446 29696 46452
rect 29736 46504 29788 46510
rect 29736 46446 29788 46452
rect 29656 46170 29684 46446
rect 29736 46368 29788 46374
rect 29736 46310 29788 46316
rect 29644 46164 29696 46170
rect 29644 46106 29696 46112
rect 29000 45960 29052 45966
rect 29000 45902 29052 45908
rect 29012 45558 29040 45902
rect 29000 45552 29052 45558
rect 29000 45494 29052 45500
rect 29748 45490 29776 46310
rect 29932 46034 29960 46990
rect 30300 46034 30328 49200
rect 33232 47048 33284 47054
rect 33232 46990 33284 46996
rect 33244 46646 33272 46990
rect 33232 46640 33284 46646
rect 33232 46582 33284 46588
rect 33520 46510 33548 49200
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 33232 46504 33284 46510
rect 33232 46446 33284 46452
rect 33508 46504 33560 46510
rect 33508 46446 33560 46452
rect 33244 46170 33272 46446
rect 35532 46368 35584 46374
rect 35532 46310 35584 46316
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 33232 46164 33284 46170
rect 33232 46106 33284 46112
rect 35544 46034 35572 46310
rect 36096 46034 36124 49200
rect 36740 46442 36768 49200
rect 37648 46504 37700 46510
rect 37648 46446 37700 46452
rect 36728 46436 36780 46442
rect 36728 46378 36780 46384
rect 29920 46028 29972 46034
rect 29920 45970 29972 45976
rect 30288 46028 30340 46034
rect 30288 45970 30340 45976
rect 35532 46028 35584 46034
rect 35532 45970 35584 45976
rect 36084 46028 36136 46034
rect 36084 45970 36136 45976
rect 29920 45892 29972 45898
rect 29920 45834 29972 45840
rect 35716 45892 35768 45898
rect 35716 45834 35768 45840
rect 29932 45626 29960 45834
rect 35728 45626 35756 45834
rect 29920 45620 29972 45626
rect 29920 45562 29972 45568
rect 35716 45620 35768 45626
rect 35716 45562 35768 45568
rect 37660 45558 37688 46446
rect 38672 46442 38700 49200
rect 39764 47048 39816 47054
rect 39764 46990 39816 46996
rect 39776 46578 39804 46990
rect 39764 46572 39816 46578
rect 39764 46514 39816 46520
rect 39948 46504 40000 46510
rect 39948 46446 40000 46452
rect 38660 46436 38712 46442
rect 38660 46378 38712 46384
rect 39960 46170 39988 46446
rect 39948 46164 40000 46170
rect 39948 46106 40000 46112
rect 40604 46034 40632 49200
rect 41892 46442 41920 49200
rect 42616 47048 42668 47054
rect 42616 46990 42668 46996
rect 44640 47048 44692 47054
rect 44640 46990 44692 46996
rect 45376 47048 45428 47054
rect 45376 46990 45428 46996
rect 42628 46578 42656 46990
rect 44652 46578 44680 46990
rect 42616 46572 42668 46578
rect 42616 46514 42668 46520
rect 44640 46572 44692 46578
rect 44640 46514 44692 46520
rect 42800 46504 42852 46510
rect 42800 46446 42852 46452
rect 41880 46436 41932 46442
rect 41880 46378 41932 46384
rect 41512 46096 41564 46102
rect 41512 46038 41564 46044
rect 40592 46028 40644 46034
rect 40592 45970 40644 45976
rect 37924 45960 37976 45966
rect 37924 45902 37976 45908
rect 40132 45960 40184 45966
rect 40132 45902 40184 45908
rect 37648 45552 37700 45558
rect 37648 45494 37700 45500
rect 37936 45490 37964 45902
rect 40144 45490 40172 45902
rect 40316 45892 40368 45898
rect 40316 45834 40368 45840
rect 29736 45484 29788 45490
rect 29736 45426 29788 45432
rect 35624 45484 35676 45490
rect 35624 45426 35676 45432
rect 36544 45484 36596 45490
rect 36544 45426 36596 45432
rect 37924 45484 37976 45490
rect 37924 45426 37976 45432
rect 40132 45484 40184 45490
rect 40132 45426 40184 45432
rect 27804 43784 27856 43790
rect 27804 43726 27856 43732
rect 27436 43716 27488 43722
rect 27436 43658 27488 43664
rect 27344 43648 27396 43654
rect 27344 43590 27396 43596
rect 27356 43314 27384 43590
rect 27344 43308 27396 43314
rect 27344 43250 27396 43256
rect 27448 43246 27476 43658
rect 29748 43382 29776 45426
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 29736 43376 29788 43382
rect 29736 43318 29788 43324
rect 28540 43308 28592 43314
rect 28540 43250 28592 43256
rect 29000 43308 29052 43314
rect 29000 43250 29052 43256
rect 30472 43308 30524 43314
rect 30472 43250 30524 43256
rect 27436 43240 27488 43246
rect 27436 43182 27488 43188
rect 27252 43104 27304 43110
rect 27252 43046 27304 43052
rect 27264 42226 27292 43046
rect 27344 42560 27396 42566
rect 27344 42502 27396 42508
rect 27252 42220 27304 42226
rect 27252 42162 27304 42168
rect 27356 41546 27384 42502
rect 27344 41540 27396 41546
rect 27344 41482 27396 41488
rect 26976 36848 27028 36854
rect 26976 36790 27028 36796
rect 26608 36712 26660 36718
rect 26608 36654 26660 36660
rect 27160 36712 27212 36718
rect 27160 36654 27212 36660
rect 26332 35284 26384 35290
rect 26332 35226 26384 35232
rect 26056 34944 26108 34950
rect 26056 34886 26108 34892
rect 25320 34740 25372 34746
rect 25320 34682 25372 34688
rect 24584 34672 24636 34678
rect 24584 34614 24636 34620
rect 24032 34604 24084 34610
rect 24032 34546 24084 34552
rect 26068 33998 26096 34886
rect 26056 33992 26108 33998
rect 26056 33934 26108 33940
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 24952 33516 25004 33522
rect 24952 33458 25004 33464
rect 24860 33312 24912 33318
rect 24860 33254 24912 33260
rect 24872 32842 24900 33254
rect 24860 32836 24912 32842
rect 24860 32778 24912 32784
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 24964 31414 24992 33458
rect 25964 33040 26016 33046
rect 25964 32982 26016 32988
rect 25976 32434 26004 32982
rect 26068 32910 26096 33934
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26068 32434 26096 32846
rect 26424 32836 26476 32842
rect 26424 32778 26476 32784
rect 26240 32768 26292 32774
rect 26240 32710 26292 32716
rect 25964 32428 26016 32434
rect 25964 32370 26016 32376
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26252 32366 26280 32710
rect 26436 32366 26464 32778
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 26424 32360 26476 32366
rect 26424 32302 26476 32308
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 24952 31408 25004 31414
rect 24952 31350 25004 31356
rect 26252 31346 26280 32166
rect 26332 31952 26384 31958
rect 26332 31894 26384 31900
rect 24308 31340 24360 31346
rect 24308 31282 24360 31288
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 23480 30388 23532 30394
rect 23480 30330 23532 30336
rect 23296 30320 23348 30326
rect 23296 30262 23348 30268
rect 23308 29646 23336 30262
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 23400 29850 23428 30194
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23492 29628 23520 30330
rect 23572 29640 23624 29646
rect 23492 29600 23572 29628
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 23308 29306 23336 29582
rect 23296 29300 23348 29306
rect 23124 29260 23296 29288
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 22664 27470 22692 28358
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22940 27674 22968 28018
rect 23020 28008 23072 28014
rect 23020 27950 23072 27956
rect 22928 27668 22980 27674
rect 22928 27610 22980 27616
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 22940 26994 22968 27610
rect 23032 27606 23060 27950
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 23124 27470 23152 29260
rect 23296 29242 23348 29248
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23400 28150 23428 28358
rect 23388 28144 23440 28150
rect 23388 28086 23440 28092
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 22940 25770 22968 26930
rect 22928 25764 22980 25770
rect 22928 25706 22980 25712
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22388 25226 22416 25638
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22940 25242 22968 25706
rect 22376 25220 22428 25226
rect 22376 25162 22428 25168
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 22388 24818 22416 25162
rect 22756 24818 22784 25230
rect 22940 25214 23060 25242
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 22940 24818 22968 25094
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 22204 23662 22232 24142
rect 22388 23730 22416 24754
rect 22756 23798 22784 24754
rect 23032 24206 23060 25214
rect 23124 24750 23152 27406
rect 23216 26926 23244 28018
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 23204 26920 23256 26926
rect 23204 26862 23256 26868
rect 23308 25294 23336 27270
rect 23400 27130 23428 28086
rect 23492 27878 23520 29600
rect 23572 29582 23624 29588
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 23952 29306 23980 29446
rect 24044 29306 24072 29582
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 24032 29300 24084 29306
rect 24032 29242 24084 29248
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23676 28762 23704 29038
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 23676 28082 23704 28562
rect 23664 28076 23716 28082
rect 23664 28018 23716 28024
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 23860 27985 23888 28018
rect 23846 27976 23902 27985
rect 23756 27940 23808 27946
rect 23846 27911 23902 27920
rect 23756 27882 23808 27888
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23388 27124 23440 27130
rect 23388 27066 23440 27072
rect 23492 26994 23520 27814
rect 23768 27538 23796 27882
rect 23572 27532 23624 27538
rect 23572 27474 23624 27480
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23584 26790 23612 27474
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23400 25498 23428 25842
rect 23940 25832 23992 25838
rect 23940 25774 23992 25780
rect 23952 25498 23980 25774
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23940 25492 23992 25498
rect 23940 25434 23992 25440
rect 24044 25294 24072 29242
rect 24122 28112 24178 28121
rect 24122 28047 24124 28056
rect 24176 28047 24178 28056
rect 24124 28018 24176 28024
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23848 25288 23900 25294
rect 23848 25230 23900 25236
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 23860 24954 23888 25230
rect 23848 24948 23900 24954
rect 23848 24890 23900 24896
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 22848 21690 22876 21966
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 23032 21570 23060 24142
rect 23124 24138 23152 24686
rect 23296 24676 23348 24682
rect 23296 24618 23348 24624
rect 23308 24274 23336 24618
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 23112 24132 23164 24138
rect 23112 24074 23164 24080
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23204 23656 23256 23662
rect 23204 23598 23256 23604
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23124 21842 23152 23462
rect 23216 23118 23244 23598
rect 23952 23186 23980 24006
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23216 22030 23244 22578
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23204 21888 23256 21894
rect 23124 21836 23204 21842
rect 23124 21830 23256 21836
rect 23124 21814 23244 21830
rect 23032 21554 23152 21570
rect 23032 21548 23164 21554
rect 23032 21542 23112 21548
rect 23112 21490 23164 21496
rect 23124 21078 23152 21490
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 23124 20466 23152 21014
rect 23216 21010 23244 21814
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 23308 20602 23336 22578
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23400 21894 23428 22374
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23400 20942 23428 21830
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23492 21554 23520 21626
rect 24044 21554 24072 25230
rect 24136 25226 24164 28018
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23492 20466 23520 21490
rect 23768 21146 23796 21490
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23860 20874 23888 21354
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5828 5234 5856 7822
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 8300 5160 8352 5166
rect 5644 5086 5764 5114
rect 8300 5102 8352 5108
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 3738 5580 4626
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5356 3664 5408 3670
rect 5644 3618 5672 4966
rect 5408 3612 5672 3618
rect 5356 3606 5672 3612
rect 5368 3590 5672 3606
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4896 2372 4948 2378
rect 4540 800 4568 2366
rect 4896 2314 4948 2320
rect 5184 800 5212 2926
rect 5644 2650 5672 3062
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5736 2582 5764 5086
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5736 2446 5764 2518
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6472 800 6500 3538
rect 6932 2378 6960 3878
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 7024 2310 7052 4558
rect 8312 4146 8340 5102
rect 10428 4146 10456 5578
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 7576 3058 7604 3878
rect 8404 3126 8432 3878
rect 10520 3602 10548 3878
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 10336 3058 10364 3470
rect 10612 3058 10640 4014
rect 12912 4010 12940 4082
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 2514 7144 2790
rect 7852 2774 7880 2926
rect 7760 2746 7880 2774
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7208 1306 7236 2450
rect 7116 1278 7236 1306
rect 7116 800 7144 1278
rect 7760 800 7788 2746
rect 10980 800 11008 3538
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2514 12480 2790
rect 12544 2582 12572 3878
rect 12912 2650 12940 3946
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3058 13032 3470
rect 13188 3126 13216 3878
rect 17420 3534 17448 5714
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20732 3534 20760 4014
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 16868 3058 16896 3470
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 3126 17080 3334
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12912 800 12940 2450
rect 13556 800 13584 2926
rect 17420 800 17448 2926
rect 19352 2446 19380 3470
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 2582 19472 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20272 2990 20300 3470
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 3126 20852 3334
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 22020 3058 22048 3470
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22204 3126 22232 3334
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19340 2440 19392 2446
rect 19720 2394 19748 2450
rect 19340 2382 19392 2388
rect 19444 2366 19748 2394
rect 19444 1306 19472 2366
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19352 1278 19472 1306
rect 19352 800 19380 1278
rect 20640 800 20668 2926
rect 22572 800 22600 2926
rect 24320 2514 24348 31282
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 26068 30394 26096 31078
rect 26056 30388 26108 30394
rect 26056 30330 26108 30336
rect 24400 30048 24452 30054
rect 24400 29990 24452 29996
rect 24412 29714 24440 29990
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24400 29708 24452 29714
rect 24400 29650 24452 29656
rect 24412 27470 24440 29650
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24596 29170 24624 29446
rect 24676 29232 24728 29238
rect 24676 29174 24728 29180
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24492 28960 24544 28966
rect 24492 28902 24544 28908
rect 24504 28558 24532 28902
rect 24596 28626 24624 29106
rect 24584 28620 24636 28626
rect 24584 28562 24636 28568
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24504 28014 24532 28494
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 24596 27606 24624 28562
rect 24688 28490 24716 29174
rect 24780 29102 24808 29718
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24676 28484 24728 28490
rect 24676 28426 24728 28432
rect 24584 27600 24636 27606
rect 24584 27542 24636 27548
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 24412 25702 24440 27406
rect 24688 26790 24716 28426
rect 24780 28121 24808 29038
rect 24952 28416 25004 28422
rect 24952 28358 25004 28364
rect 24964 28150 24992 28358
rect 26344 28150 26372 31894
rect 26516 31816 26568 31822
rect 26516 31758 26568 31764
rect 26528 31346 26556 31758
rect 26620 31754 26648 36654
rect 27172 36038 27200 36654
rect 27344 36576 27396 36582
rect 27344 36518 27396 36524
rect 27160 36032 27212 36038
rect 27160 35974 27212 35980
rect 27356 35698 27384 36518
rect 27344 35692 27396 35698
rect 27344 35634 27396 35640
rect 26700 35284 26752 35290
rect 26700 35226 26752 35232
rect 26712 33454 26740 35226
rect 27448 34610 27476 43182
rect 28552 42770 28580 43250
rect 28080 42764 28132 42770
rect 28080 42706 28132 42712
rect 28540 42764 28592 42770
rect 28540 42706 28592 42712
rect 28092 42294 28120 42706
rect 28448 42696 28500 42702
rect 28448 42638 28500 42644
rect 28724 42696 28776 42702
rect 28724 42638 28776 42644
rect 28080 42288 28132 42294
rect 28080 42230 28132 42236
rect 27896 42016 27948 42022
rect 27896 41958 27948 41964
rect 27908 41414 27936 41958
rect 28092 41614 28120 42230
rect 28460 41818 28488 42638
rect 28736 42294 28764 42638
rect 28908 42628 28960 42634
rect 28908 42570 28960 42576
rect 28724 42288 28776 42294
rect 28724 42230 28776 42236
rect 28540 42016 28592 42022
rect 28540 41958 28592 41964
rect 28448 41812 28500 41818
rect 28448 41754 28500 41760
rect 28080 41608 28132 41614
rect 28080 41550 28132 41556
rect 27908 41386 28028 41414
rect 27804 39296 27856 39302
rect 27804 39238 27856 39244
rect 27816 38350 27844 39238
rect 27804 38344 27856 38350
rect 27804 38286 27856 38292
rect 28000 37330 28028 41386
rect 28092 39982 28120 41550
rect 28552 40730 28580 41958
rect 28632 41812 28684 41818
rect 28632 41754 28684 41760
rect 28264 40724 28316 40730
rect 28264 40666 28316 40672
rect 28540 40724 28592 40730
rect 28540 40666 28592 40672
rect 28080 39976 28132 39982
rect 28080 39918 28132 39924
rect 28092 38962 28120 39918
rect 28276 39506 28304 40666
rect 28644 40662 28672 41754
rect 28736 41614 28764 42230
rect 28920 41818 28948 42570
rect 29012 42090 29040 43250
rect 29828 43104 29880 43110
rect 29828 43046 29880 43052
rect 30288 43104 30340 43110
rect 30288 43046 30340 43052
rect 29184 42560 29236 42566
rect 29184 42502 29236 42508
rect 29196 42226 29224 42502
rect 29840 42226 29868 43046
rect 30300 42702 30328 43046
rect 30288 42696 30340 42702
rect 30288 42638 30340 42644
rect 30484 42294 30512 43250
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 32128 42696 32180 42702
rect 32128 42638 32180 42644
rect 35348 42696 35400 42702
rect 35348 42638 35400 42644
rect 31116 42560 31168 42566
rect 31116 42502 31168 42508
rect 30472 42288 30524 42294
rect 30472 42230 30524 42236
rect 31128 42226 31156 42502
rect 29184 42220 29236 42226
rect 29184 42162 29236 42168
rect 29828 42220 29880 42226
rect 29828 42162 29880 42168
rect 31116 42220 31168 42226
rect 31116 42162 31168 42168
rect 30564 42152 30616 42158
rect 30564 42094 30616 42100
rect 29000 42084 29052 42090
rect 29000 42026 29052 42032
rect 28908 41812 28960 41818
rect 28908 41754 28960 41760
rect 30576 41614 30604 42094
rect 31128 41750 31156 42162
rect 31116 41744 31168 41750
rect 31116 41686 31168 41692
rect 28724 41608 28776 41614
rect 28724 41550 28776 41556
rect 30564 41608 30616 41614
rect 30564 41550 30616 41556
rect 29920 41540 29972 41546
rect 29920 41482 29972 41488
rect 29932 40730 29960 41482
rect 30576 40934 30604 41550
rect 30656 41540 30708 41546
rect 30656 41482 30708 41488
rect 31024 41540 31076 41546
rect 31024 41482 31076 41488
rect 30668 41070 30696 41482
rect 30932 41472 30984 41478
rect 30932 41414 30984 41420
rect 30944 41206 30972 41414
rect 30932 41200 30984 41206
rect 30932 41142 30984 41148
rect 30656 41064 30708 41070
rect 30656 41006 30708 41012
rect 30564 40928 30616 40934
rect 30564 40870 30616 40876
rect 30840 40928 30892 40934
rect 30840 40870 30892 40876
rect 29920 40724 29972 40730
rect 29920 40666 29972 40672
rect 28632 40656 28684 40662
rect 28632 40598 28684 40604
rect 28264 39500 28316 39506
rect 28264 39442 28316 39448
rect 28644 39438 28672 40598
rect 29736 40452 29788 40458
rect 29736 40394 29788 40400
rect 29748 39438 29776 40394
rect 29828 40384 29880 40390
rect 29828 40326 29880 40332
rect 29840 39982 29868 40326
rect 29932 40186 29960 40666
rect 30104 40384 30156 40390
rect 30104 40326 30156 40332
rect 29920 40180 29972 40186
rect 29920 40122 29972 40128
rect 30012 40044 30064 40050
rect 30012 39986 30064 39992
rect 29828 39976 29880 39982
rect 29828 39918 29880 39924
rect 30024 39642 30052 39986
rect 30012 39636 30064 39642
rect 30012 39578 30064 39584
rect 30116 39506 30144 40326
rect 30852 40050 30880 40870
rect 31036 40458 31064 41482
rect 31128 41138 31156 41686
rect 31484 41676 31536 41682
rect 31484 41618 31536 41624
rect 31116 41132 31168 41138
rect 31116 41074 31168 41080
rect 31024 40452 31076 40458
rect 31024 40394 31076 40400
rect 30840 40044 30892 40050
rect 30840 39986 30892 39992
rect 30932 40044 30984 40050
rect 30932 39986 30984 39992
rect 30380 39908 30432 39914
rect 30380 39850 30432 39856
rect 30104 39500 30156 39506
rect 30104 39442 30156 39448
rect 30392 39438 30420 39850
rect 30472 39840 30524 39846
rect 30472 39782 30524 39788
rect 28172 39432 28224 39438
rect 28172 39374 28224 39380
rect 28632 39432 28684 39438
rect 28632 39374 28684 39380
rect 28908 39432 28960 39438
rect 28908 39374 28960 39380
rect 29736 39432 29788 39438
rect 29736 39374 29788 39380
rect 30380 39432 30432 39438
rect 30380 39374 30432 39380
rect 28080 38956 28132 38962
rect 28080 38898 28132 38904
rect 28092 37874 28120 38898
rect 28080 37868 28132 37874
rect 28080 37810 28132 37816
rect 27528 37324 27580 37330
rect 27528 37266 27580 37272
rect 27988 37324 28040 37330
rect 27988 37266 28040 37272
rect 27540 35834 27568 37266
rect 27528 35828 27580 35834
rect 27528 35770 27580 35776
rect 28000 35494 28028 37266
rect 28092 35698 28120 37810
rect 28184 37262 28212 39374
rect 28540 39364 28592 39370
rect 28540 39306 28592 39312
rect 28356 39296 28408 39302
rect 28356 39238 28408 39244
rect 28368 37874 28396 39238
rect 28552 39030 28580 39306
rect 28920 39030 28948 39374
rect 29748 39098 29776 39374
rect 30484 39370 30512 39782
rect 30472 39364 30524 39370
rect 30472 39306 30524 39312
rect 29736 39092 29788 39098
rect 29736 39034 29788 39040
rect 28540 39024 28592 39030
rect 28540 38966 28592 38972
rect 28908 39024 28960 39030
rect 28908 38966 28960 38972
rect 28552 38554 28580 38966
rect 28540 38548 28592 38554
rect 28540 38490 28592 38496
rect 28356 37868 28408 37874
rect 28356 37810 28408 37816
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 28184 36922 28212 37198
rect 28920 37194 28948 38966
rect 30944 38010 30972 39986
rect 31496 39438 31524 41618
rect 32140 41614 32168 42638
rect 32864 42628 32916 42634
rect 32864 42570 32916 42576
rect 33876 42628 33928 42634
rect 33876 42570 33928 42576
rect 32404 42560 32456 42566
rect 32404 42502 32456 42508
rect 32312 42016 32364 42022
rect 32312 41958 32364 41964
rect 32128 41608 32180 41614
rect 32128 41550 32180 41556
rect 32140 40594 32168 41550
rect 32324 41546 32352 41958
rect 32312 41540 32364 41546
rect 32312 41482 32364 41488
rect 32416 41138 32444 42502
rect 32876 42362 32904 42570
rect 32864 42356 32916 42362
rect 32864 42298 32916 42304
rect 33888 42226 33916 42570
rect 34888 42560 34940 42566
rect 34888 42502 34940 42508
rect 34900 42226 34928 42502
rect 32496 42220 32548 42226
rect 32496 42162 32548 42168
rect 33876 42220 33928 42226
rect 33876 42162 33928 42168
rect 34888 42220 34940 42226
rect 34888 42162 34940 42168
rect 32508 41274 32536 42162
rect 33140 42084 33192 42090
rect 33140 42026 33192 42032
rect 33152 41274 33180 42026
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41818 35388 42638
rect 35532 42016 35584 42022
rect 35532 41958 35584 41964
rect 35348 41812 35400 41818
rect 35348 41754 35400 41760
rect 34796 41608 34848 41614
rect 34796 41550 34848 41556
rect 34060 41540 34112 41546
rect 34060 41482 34112 41488
rect 34072 41274 34100 41482
rect 32496 41268 32548 41274
rect 32496 41210 32548 41216
rect 33140 41268 33192 41274
rect 33140 41210 33192 41216
rect 34060 41268 34112 41274
rect 34060 41210 34112 41216
rect 32404 41132 32456 41138
rect 32404 41074 32456 41080
rect 33968 41132 34020 41138
rect 33968 41074 34020 41080
rect 33784 40928 33836 40934
rect 33784 40870 33836 40876
rect 32128 40588 32180 40594
rect 32128 40530 32180 40536
rect 32956 40588 33008 40594
rect 32956 40530 33008 40536
rect 31300 39432 31352 39438
rect 31300 39374 31352 39380
rect 31484 39432 31536 39438
rect 31484 39374 31536 39380
rect 32036 39432 32088 39438
rect 32036 39374 32088 39380
rect 31208 38956 31260 38962
rect 31208 38898 31260 38904
rect 31116 38752 31168 38758
rect 31116 38694 31168 38700
rect 31128 38350 31156 38694
rect 31116 38344 31168 38350
rect 31116 38286 31168 38292
rect 31220 38010 31248 38898
rect 31312 38758 31340 39374
rect 32048 38962 32076 39374
rect 32036 38956 32088 38962
rect 32036 38898 32088 38904
rect 31300 38752 31352 38758
rect 31300 38694 31352 38700
rect 29460 38004 29512 38010
rect 29460 37946 29512 37952
rect 30932 38004 30984 38010
rect 30932 37946 30984 37952
rect 31208 38004 31260 38010
rect 31208 37946 31260 37952
rect 28908 37188 28960 37194
rect 28908 37130 28960 37136
rect 28448 37120 28500 37126
rect 28448 37062 28500 37068
rect 28172 36916 28224 36922
rect 28172 36858 28224 36864
rect 28264 36780 28316 36786
rect 28264 36722 28316 36728
rect 28276 36378 28304 36722
rect 28264 36372 28316 36378
rect 28264 36314 28316 36320
rect 28460 36174 28488 37062
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 28080 35692 28132 35698
rect 28080 35634 28132 35640
rect 29276 35692 29328 35698
rect 29276 35634 29328 35640
rect 27988 35488 28040 35494
rect 27988 35430 28040 35436
rect 27528 34672 27580 34678
rect 27528 34614 27580 34620
rect 27436 34604 27488 34610
rect 27436 34546 27488 34552
rect 27344 34400 27396 34406
rect 27344 34342 27396 34348
rect 27160 33924 27212 33930
rect 27160 33866 27212 33872
rect 27068 33856 27120 33862
rect 27068 33798 27120 33804
rect 26700 33448 26752 33454
rect 26700 33390 26752 33396
rect 26712 33046 26740 33390
rect 26700 33040 26752 33046
rect 26700 32982 26752 32988
rect 26712 32366 26740 32982
rect 26884 32768 26936 32774
rect 26884 32710 26936 32716
rect 26700 32360 26752 32366
rect 26700 32302 26752 32308
rect 26792 32224 26844 32230
rect 26792 32166 26844 32172
rect 26804 31754 26832 32166
rect 26620 31726 26740 31754
rect 26608 31680 26660 31686
rect 26608 31622 26660 31628
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26528 30734 26556 31282
rect 26620 31278 26648 31622
rect 26608 31272 26660 31278
rect 26608 31214 26660 31220
rect 26620 30734 26648 31214
rect 26516 30728 26568 30734
rect 26516 30670 26568 30676
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26608 30592 26660 30598
rect 26608 30534 26660 30540
rect 26620 29646 26648 30534
rect 26608 29640 26660 29646
rect 26608 29582 26660 29588
rect 26424 29572 26476 29578
rect 26424 29514 26476 29520
rect 26436 29170 26464 29514
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26528 28558 26556 29446
rect 26608 29164 26660 29170
rect 26608 29106 26660 29112
rect 26620 28762 26648 29106
rect 26608 28756 26660 28762
rect 26608 28698 26660 28704
rect 26712 28694 26740 31726
rect 26792 31748 26844 31754
rect 26792 31690 26844 31696
rect 26804 30734 26832 31690
rect 26896 31686 26924 32710
rect 27080 32570 27108 33798
rect 27172 33658 27200 33866
rect 27160 33652 27212 33658
rect 27160 33594 27212 33600
rect 27356 33522 27384 34342
rect 27448 33590 27476 34546
rect 27436 33584 27488 33590
rect 27436 33526 27488 33532
rect 27344 33516 27396 33522
rect 27344 33458 27396 33464
rect 27540 32842 27568 34614
rect 28092 34610 28120 35634
rect 29288 35290 29316 35634
rect 29276 35284 29328 35290
rect 29276 35226 29328 35232
rect 29472 34678 29500 37946
rect 31208 37868 31260 37874
rect 31312 37856 31340 38694
rect 31260 37828 31340 37856
rect 31208 37810 31260 37816
rect 31024 37800 31076 37806
rect 31024 37742 31076 37748
rect 31036 37466 31064 37742
rect 31024 37460 31076 37466
rect 31024 37402 31076 37408
rect 31220 36786 31248 37810
rect 32048 36854 32076 38898
rect 32140 38554 32168 40530
rect 32968 40050 32996 40530
rect 33796 40526 33824 40870
rect 33784 40520 33836 40526
rect 33784 40462 33836 40468
rect 32956 40044 33008 40050
rect 33232 40044 33284 40050
rect 33008 40004 33088 40032
rect 32956 39986 33008 39992
rect 33060 38894 33088 40004
rect 33232 39986 33284 39992
rect 33244 39642 33272 39986
rect 33980 39642 34008 41074
rect 33232 39636 33284 39642
rect 33232 39578 33284 39584
rect 33968 39636 34020 39642
rect 33968 39578 34020 39584
rect 34072 39438 34100 41210
rect 34808 40730 34836 41550
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34796 40724 34848 40730
rect 34796 40666 34848 40672
rect 34520 40452 34572 40458
rect 34520 40394 34572 40400
rect 34532 40186 34560 40394
rect 35348 40384 35400 40390
rect 35348 40326 35400 40332
rect 34520 40180 34572 40186
rect 34520 40122 34572 40128
rect 34060 39432 34112 39438
rect 34060 39374 34112 39380
rect 34072 39302 34100 39374
rect 34532 39370 34560 40122
rect 35360 40118 35388 40326
rect 35544 40118 35572 41958
rect 35636 41274 35664 45426
rect 36084 43308 36136 43314
rect 36084 43250 36136 43256
rect 35900 43104 35952 43110
rect 35900 43046 35952 43052
rect 35912 42702 35940 43046
rect 35900 42696 35952 42702
rect 35900 42638 35952 42644
rect 36096 42362 36124 43250
rect 36084 42356 36136 42362
rect 36084 42298 36136 42304
rect 36556 42294 36584 45426
rect 40328 45082 40356 45834
rect 41524 45490 41552 46038
rect 42812 45558 42840 46446
rect 45388 46102 45416 46990
rect 45560 46980 45612 46986
rect 45560 46922 45612 46928
rect 45572 46170 45600 46922
rect 45744 46368 45796 46374
rect 45744 46310 45796 46316
rect 45560 46164 45612 46170
rect 45560 46106 45612 46112
rect 45376 46096 45428 46102
rect 45376 46038 45428 46044
rect 45756 46034 45784 46310
rect 45744 46028 45796 46034
rect 45744 45970 45796 45976
rect 42800 45552 42852 45558
rect 45848 45554 45876 49286
rect 46358 49200 46470 49286
rect 47002 49200 47114 49800
rect 48290 49200 48402 49800
rect 48934 49200 49046 49800
rect 49578 49200 49690 49800
rect 46846 46336 46902 46345
rect 46846 46271 46902 46280
rect 45928 45892 45980 45898
rect 45928 45834 45980 45840
rect 42800 45494 42852 45500
rect 45756 45526 45876 45554
rect 41512 45484 41564 45490
rect 41512 45426 41564 45432
rect 40316 45076 40368 45082
rect 40316 45018 40368 45024
rect 40224 44872 40276 44878
rect 40224 44814 40276 44820
rect 40236 44334 40264 44814
rect 41524 44402 41552 45426
rect 41512 44396 41564 44402
rect 41512 44338 41564 44344
rect 40224 44328 40276 44334
rect 40224 44270 40276 44276
rect 37188 42560 37240 42566
rect 37188 42502 37240 42508
rect 36544 42288 36596 42294
rect 36544 42230 36596 42236
rect 35900 42220 35952 42226
rect 35900 42162 35952 42168
rect 35912 41818 35940 42162
rect 37200 42158 37228 42502
rect 37648 42220 37700 42226
rect 37648 42162 37700 42168
rect 38568 42220 38620 42226
rect 38568 42162 38620 42168
rect 43444 42220 43496 42226
rect 43444 42162 43496 42168
rect 37188 42152 37240 42158
rect 37188 42094 37240 42100
rect 36728 42016 36780 42022
rect 36728 41958 36780 41964
rect 35900 41812 35952 41818
rect 35900 41754 35952 41760
rect 36740 41546 36768 41958
rect 36728 41540 36780 41546
rect 36728 41482 36780 41488
rect 35624 41268 35676 41274
rect 35624 41210 35676 41216
rect 36544 41064 36596 41070
rect 36544 41006 36596 41012
rect 35808 40724 35860 40730
rect 35808 40666 35860 40672
rect 35820 40186 35848 40666
rect 36556 40390 36584 41006
rect 37200 41002 37228 42094
rect 37660 41818 37688 42162
rect 38292 42016 38344 42022
rect 38292 41958 38344 41964
rect 37648 41812 37700 41818
rect 37648 41754 37700 41760
rect 37660 41614 37688 41754
rect 38200 41676 38252 41682
rect 38200 41618 38252 41624
rect 37464 41608 37516 41614
rect 37464 41550 37516 41556
rect 37648 41608 37700 41614
rect 37648 41550 37700 41556
rect 37372 41200 37424 41206
rect 37372 41142 37424 41148
rect 37280 41132 37332 41138
rect 37280 41074 37332 41080
rect 37188 40996 37240 41002
rect 37188 40938 37240 40944
rect 36636 40928 36688 40934
rect 37200 40882 37228 40938
rect 36636 40870 36688 40876
rect 36544 40384 36596 40390
rect 36544 40326 36596 40332
rect 35808 40180 35860 40186
rect 35808 40122 35860 40128
rect 35348 40112 35400 40118
rect 35348 40054 35400 40060
rect 35532 40112 35584 40118
rect 35532 40054 35584 40060
rect 35440 39908 35492 39914
rect 35440 39850 35492 39856
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35452 39642 35480 39850
rect 35440 39636 35492 39642
rect 35440 39578 35492 39584
rect 35544 39506 35572 40054
rect 36648 40050 36676 40870
rect 37108 40854 37228 40882
rect 37108 40458 37136 40854
rect 37292 40662 37320 41074
rect 37384 41070 37412 41142
rect 37476 41070 37504 41550
rect 38212 41478 38240 41618
rect 37740 41472 37792 41478
rect 37740 41414 37792 41420
rect 38200 41472 38252 41478
rect 38200 41414 38252 41420
rect 37752 41138 37780 41414
rect 38304 41206 38332 41958
rect 38580 41818 38608 42162
rect 38752 42152 38804 42158
rect 38752 42094 38804 42100
rect 42616 42152 42668 42158
rect 42616 42094 42668 42100
rect 38568 41812 38620 41818
rect 38568 41754 38620 41760
rect 38292 41200 38344 41206
rect 38292 41142 38344 41148
rect 37740 41132 37792 41138
rect 37740 41074 37792 41080
rect 37372 41064 37424 41070
rect 37372 41006 37424 41012
rect 37464 41064 37516 41070
rect 37464 41006 37516 41012
rect 37280 40656 37332 40662
rect 37280 40598 37332 40604
rect 37384 40458 37412 41006
rect 38568 40928 38620 40934
rect 38568 40870 38620 40876
rect 38580 40594 38608 40870
rect 38568 40588 38620 40594
rect 38568 40530 38620 40536
rect 37096 40452 37148 40458
rect 37096 40394 37148 40400
rect 37372 40452 37424 40458
rect 37372 40394 37424 40400
rect 37188 40384 37240 40390
rect 37188 40326 37240 40332
rect 37200 40186 37228 40326
rect 37188 40180 37240 40186
rect 37188 40122 37240 40128
rect 36636 40044 36688 40050
rect 36636 39986 36688 39992
rect 36728 40044 36780 40050
rect 36728 39986 36780 39992
rect 35808 39976 35860 39982
rect 35808 39918 35860 39924
rect 35716 39840 35768 39846
rect 35716 39782 35768 39788
rect 35532 39500 35584 39506
rect 35532 39442 35584 39448
rect 34520 39364 34572 39370
rect 34520 39306 34572 39312
rect 34060 39296 34112 39302
rect 34060 39238 34112 39244
rect 35728 39030 35756 39782
rect 35716 39024 35768 39030
rect 35716 38966 35768 38972
rect 33048 38888 33100 38894
rect 33048 38830 33100 38836
rect 34612 38820 34664 38826
rect 34612 38762 34664 38768
rect 32864 38752 32916 38758
rect 32864 38694 32916 38700
rect 32128 38548 32180 38554
rect 32128 38490 32180 38496
rect 32140 37874 32168 38490
rect 32876 38350 32904 38694
rect 33416 38412 33468 38418
rect 33416 38354 33468 38360
rect 32864 38344 32916 38350
rect 32864 38286 32916 38292
rect 32128 37868 32180 37874
rect 32128 37810 32180 37816
rect 32140 37262 32168 37810
rect 33048 37392 33100 37398
rect 33048 37334 33100 37340
rect 32128 37256 32180 37262
rect 32128 37198 32180 37204
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32140 36854 32168 37198
rect 32324 36922 32352 37198
rect 32312 36916 32364 36922
rect 32312 36858 32364 36864
rect 32036 36848 32088 36854
rect 32036 36790 32088 36796
rect 32128 36848 32180 36854
rect 32128 36790 32180 36796
rect 30656 36780 30708 36786
rect 30656 36722 30708 36728
rect 31208 36780 31260 36786
rect 31208 36722 31260 36728
rect 30564 35488 30616 35494
rect 30564 35430 30616 35436
rect 30576 35154 30604 35430
rect 30564 35148 30616 35154
rect 30564 35090 30616 35096
rect 30472 35080 30524 35086
rect 30472 35022 30524 35028
rect 30380 35012 30432 35018
rect 30380 34954 30432 34960
rect 30392 34746 30420 34954
rect 30380 34740 30432 34746
rect 30380 34682 30432 34688
rect 29460 34672 29512 34678
rect 29460 34614 29512 34620
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 28920 34202 28948 34546
rect 28908 34196 28960 34202
rect 28908 34138 28960 34144
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 30380 33992 30432 33998
rect 30484 33980 30512 35022
rect 30576 33998 30604 35090
rect 30432 33952 30512 33980
rect 30564 33992 30616 33998
rect 30380 33934 30432 33940
rect 30564 33934 30616 33940
rect 29840 33522 29868 33934
rect 29828 33516 29880 33522
rect 29828 33458 29880 33464
rect 27528 32836 27580 32842
rect 27528 32778 27580 32784
rect 27068 32564 27120 32570
rect 27068 32506 27120 32512
rect 27080 31822 27108 32506
rect 27540 32298 27568 32778
rect 29736 32768 29788 32774
rect 29736 32710 29788 32716
rect 29748 32502 29776 32710
rect 29840 32570 29868 33458
rect 29828 32564 29880 32570
rect 29828 32506 29880 32512
rect 29736 32496 29788 32502
rect 29736 32438 29788 32444
rect 27252 32292 27304 32298
rect 27252 32234 27304 32240
rect 27528 32292 27580 32298
rect 27528 32234 27580 32240
rect 27264 31822 27292 32234
rect 27620 32224 27672 32230
rect 27620 32166 27672 32172
rect 27068 31816 27120 31822
rect 27068 31758 27120 31764
rect 27252 31816 27304 31822
rect 27252 31758 27304 31764
rect 26976 31748 27028 31754
rect 26976 31690 27028 31696
rect 26884 31680 26936 31686
rect 26884 31622 26936 31628
rect 26988 31482 27016 31690
rect 27528 31680 27580 31686
rect 27528 31622 27580 31628
rect 26976 31476 27028 31482
rect 26976 31418 27028 31424
rect 27540 31414 27568 31622
rect 27528 31408 27580 31414
rect 27528 31350 27580 31356
rect 27632 31346 27660 32166
rect 30392 31822 30420 33934
rect 30576 33590 30604 33934
rect 30564 33584 30616 33590
rect 30564 33526 30616 33532
rect 30564 32904 30616 32910
rect 30564 32846 30616 32852
rect 30576 32026 30604 32846
rect 30564 32020 30616 32026
rect 30564 31962 30616 31968
rect 29092 31816 29144 31822
rect 29092 31758 29144 31764
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27172 30734 27200 31282
rect 29104 31278 29132 31758
rect 29736 31680 29788 31686
rect 29736 31622 29788 31628
rect 29748 31482 29776 31622
rect 29736 31476 29788 31482
rect 29736 31418 29788 31424
rect 29092 31272 29144 31278
rect 29092 31214 29144 31220
rect 29368 31272 29420 31278
rect 29368 31214 29420 31220
rect 27896 31136 27948 31142
rect 27896 31078 27948 31084
rect 26792 30728 26844 30734
rect 26792 30670 26844 30676
rect 27160 30728 27212 30734
rect 27160 30670 27212 30676
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27448 29850 27476 30670
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27160 29572 27212 29578
rect 27160 29514 27212 29520
rect 27172 29306 27200 29514
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 27448 29170 27476 29786
rect 27908 29510 27936 31078
rect 28724 29640 28776 29646
rect 28724 29582 28776 29588
rect 27896 29504 27948 29510
rect 27896 29446 27948 29452
rect 28736 29170 28764 29582
rect 29380 29238 29408 31214
rect 29748 30802 29776 31418
rect 30208 31414 30236 31758
rect 30196 31408 30248 31414
rect 30196 31350 30248 31356
rect 30104 31340 30156 31346
rect 30104 31282 30156 31288
rect 30116 30938 30144 31282
rect 30104 30932 30156 30938
rect 30104 30874 30156 30880
rect 29736 30796 29788 30802
rect 29736 30738 29788 30744
rect 30392 30734 30420 31758
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30012 30388 30064 30394
rect 30012 30330 30064 30336
rect 29368 29232 29420 29238
rect 29368 29174 29420 29180
rect 29828 29232 29880 29238
rect 29828 29174 29880 29180
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27620 29164 27672 29170
rect 27620 29106 27672 29112
rect 28724 29164 28776 29170
rect 28724 29106 28776 29112
rect 26792 28960 26844 28966
rect 26792 28902 26844 28908
rect 26700 28688 26752 28694
rect 26700 28630 26752 28636
rect 26804 28626 26832 28902
rect 26792 28620 26844 28626
rect 26792 28562 26844 28568
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 24952 28144 25004 28150
rect 24766 28112 24822 28121
rect 24952 28086 25004 28092
rect 25596 28144 25648 28150
rect 25596 28086 25648 28092
rect 26332 28144 26384 28150
rect 26332 28086 26384 28092
rect 24766 28047 24822 28056
rect 25226 27976 25282 27985
rect 24768 27940 24820 27946
rect 25226 27911 25228 27920
rect 24768 27882 24820 27888
rect 25280 27911 25282 27920
rect 25228 27882 25280 27888
rect 24780 26926 24808 27882
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24872 27470 24900 27814
rect 25608 27606 25636 28086
rect 25596 27600 25648 27606
rect 25596 27542 25648 27548
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 25608 27402 25636 27542
rect 26344 27538 26372 28086
rect 26528 28082 26556 28494
rect 27448 28490 27476 29106
rect 27632 28762 27660 29106
rect 27896 28960 27948 28966
rect 27896 28902 27948 28908
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 27908 28558 27936 28902
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 27436 28484 27488 28490
rect 27436 28426 27488 28432
rect 26608 28416 26660 28422
rect 26608 28358 26660 28364
rect 26620 28150 26648 28358
rect 26608 28144 26660 28150
rect 26608 28086 26660 28092
rect 26516 28076 26568 28082
rect 26516 28018 26568 28024
rect 26620 27674 26648 28086
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 26332 27532 26384 27538
rect 26332 27474 26384 27480
rect 25596 27396 25648 27402
rect 25596 27338 25648 27344
rect 25688 27396 25740 27402
rect 25688 27338 25740 27344
rect 25700 27062 25728 27338
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25688 27056 25740 27062
rect 25688 26998 25740 27004
rect 25976 26994 26004 27270
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 26344 26926 26372 27474
rect 26608 27464 26660 27470
rect 27448 27452 27476 28426
rect 28540 27872 28592 27878
rect 28540 27814 28592 27820
rect 27528 27464 27580 27470
rect 27448 27424 27528 27452
rect 26608 27406 26660 27412
rect 27528 27406 27580 27412
rect 26620 27130 26648 27406
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 26608 27124 26660 27130
rect 26608 27066 26660 27072
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27528 26988 27580 26994
rect 27632 26976 27660 27270
rect 27580 26948 27660 26976
rect 27528 26930 27580 26936
rect 24768 26920 24820 26926
rect 24768 26862 24820 26868
rect 26332 26920 26384 26926
rect 27448 26897 27476 26930
rect 26332 26862 26384 26868
rect 27434 26888 27490 26897
rect 27344 26852 27396 26858
rect 27434 26823 27490 26832
rect 27344 26794 27396 26800
rect 24676 26784 24728 26790
rect 24676 26726 24728 26732
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 26344 25838 26372 26318
rect 27356 26246 27384 26794
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 27448 26382 27476 26726
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27344 26240 27396 26246
rect 27344 26182 27396 26188
rect 27356 25906 27384 26182
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 26332 25832 26384 25838
rect 27632 25820 27660 26948
rect 27804 26988 27856 26994
rect 27804 26930 27856 26936
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 27724 26382 27752 26726
rect 27816 26382 27844 26930
rect 27894 26888 27950 26897
rect 27894 26823 27950 26832
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27804 26376 27856 26382
rect 27804 26318 27856 26324
rect 27804 26240 27856 26246
rect 27804 26182 27856 26188
rect 27816 25974 27844 26182
rect 27804 25968 27856 25974
rect 27804 25910 27856 25916
rect 27632 25792 27844 25820
rect 26332 25774 26384 25780
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 24412 23118 24440 25638
rect 25424 25294 25452 25638
rect 26344 25498 26372 25774
rect 27436 25696 27488 25702
rect 27436 25638 27488 25644
rect 27712 25696 27764 25702
rect 27712 25638 27764 25644
rect 26332 25492 26384 25498
rect 26332 25434 26384 25440
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 24964 24410 24992 25230
rect 25320 25220 25372 25226
rect 25320 25162 25372 25168
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24596 23730 24624 24006
rect 25332 23730 25360 25162
rect 27448 24750 27476 25638
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 27632 24818 27660 25094
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27436 24744 27488 24750
rect 27436 24686 27488 24692
rect 27448 24206 27476 24686
rect 27724 24342 27752 25638
rect 27816 25226 27844 25792
rect 27908 25294 27936 26823
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 27804 25220 27856 25226
rect 27804 25162 27856 25168
rect 27908 24954 27936 25230
rect 27896 24948 27948 24954
rect 27896 24890 27948 24896
rect 27804 24812 27856 24818
rect 27804 24754 27856 24760
rect 27896 24812 27948 24818
rect 27896 24754 27948 24760
rect 27816 24410 27844 24754
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27712 24336 27764 24342
rect 27712 24278 27764 24284
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 27252 24200 27304 24206
rect 27252 24142 27304 24148
rect 27436 24200 27488 24206
rect 27436 24142 27488 24148
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25516 23730 25544 24006
rect 26160 23730 26188 24142
rect 26884 24132 26936 24138
rect 26884 24074 26936 24080
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 24872 23322 24900 23666
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24964 23118 24992 23462
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24412 21554 24440 23054
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24412 21078 24440 21490
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 25332 20874 25360 23666
rect 26160 23322 26188 23666
rect 26148 23316 26200 23322
rect 26148 23258 26200 23264
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 26240 22092 26292 22098
rect 26240 22034 26292 22040
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 26252 20466 26280 22034
rect 26436 21690 26464 22578
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 26896 21554 26924 24074
rect 27264 23866 27292 24142
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 26976 23656 27028 23662
rect 26976 23598 27028 23604
rect 26988 23118 27016 23598
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 26988 22234 27016 23054
rect 27080 22778 27108 23054
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 27540 22658 27568 24074
rect 27632 22778 27660 24142
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27724 23186 27752 23598
rect 27816 23254 27844 24006
rect 27908 23322 27936 24754
rect 28000 23866 28028 25842
rect 28092 25498 28120 26386
rect 28080 25492 28132 25498
rect 28080 25434 28132 25440
rect 28184 25362 28212 27270
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28080 25152 28132 25158
rect 28080 25094 28132 25100
rect 28092 24682 28120 25094
rect 28184 24818 28212 25298
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28080 24676 28132 24682
rect 28080 24618 28132 24624
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 28092 23526 28120 24618
rect 28552 24206 28580 27814
rect 29840 27538 29868 29174
rect 29920 29096 29972 29102
rect 29920 29038 29972 29044
rect 29932 28966 29960 29038
rect 29920 28960 29972 28966
rect 29920 28902 29972 28908
rect 29932 28422 29960 28902
rect 30024 28558 30052 30330
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 30668 28490 30696 36722
rect 32140 36378 32168 36790
rect 33060 36718 33088 37334
rect 33324 37256 33376 37262
rect 33324 37198 33376 37204
rect 33140 37188 33192 37194
rect 33140 37130 33192 37136
rect 33152 36786 33180 37130
rect 33232 37120 33284 37126
rect 33232 37062 33284 37068
rect 33140 36780 33192 36786
rect 33140 36722 33192 36728
rect 33048 36712 33100 36718
rect 33048 36654 33100 36660
rect 33244 36582 33272 37062
rect 33336 36786 33364 37198
rect 33428 37194 33456 38354
rect 33508 38208 33560 38214
rect 33508 38150 33560 38156
rect 33520 37942 33548 38150
rect 33508 37936 33560 37942
rect 33508 37878 33560 37884
rect 33968 37664 34020 37670
rect 33968 37606 34020 37612
rect 33980 37262 34008 37606
rect 34624 37398 34652 38762
rect 35820 38758 35848 39918
rect 36740 39098 36768 39986
rect 38580 39982 38608 40530
rect 38108 39976 38160 39982
rect 38108 39918 38160 39924
rect 38568 39976 38620 39982
rect 38568 39918 38620 39924
rect 38120 39438 38148 39918
rect 38108 39432 38160 39438
rect 38108 39374 38160 39380
rect 37556 39364 37608 39370
rect 37556 39306 37608 39312
rect 36728 39092 36780 39098
rect 36728 39034 36780 39040
rect 35808 38752 35860 38758
rect 35808 38694 35860 38700
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 36740 38418 36768 39034
rect 37568 38962 37596 39306
rect 37556 38956 37608 38962
rect 37556 38898 37608 38904
rect 36728 38412 36780 38418
rect 36728 38354 36780 38360
rect 37188 38412 37240 38418
rect 37188 38354 37240 38360
rect 37096 38344 37148 38350
rect 37096 38286 37148 38292
rect 36912 38208 36964 38214
rect 36912 38150 36964 38156
rect 36924 37874 36952 38150
rect 36912 37868 36964 37874
rect 36912 37810 36964 37816
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35440 37460 35492 37466
rect 35440 37402 35492 37408
rect 34612 37392 34664 37398
rect 34612 37334 34664 37340
rect 34704 37324 34756 37330
rect 34704 37266 34756 37272
rect 33968 37256 34020 37262
rect 33968 37198 34020 37204
rect 33416 37188 33468 37194
rect 33416 37130 33468 37136
rect 33324 36780 33376 36786
rect 33324 36722 33376 36728
rect 33140 36576 33192 36582
rect 33140 36518 33192 36524
rect 33232 36576 33284 36582
rect 33232 36518 33284 36524
rect 33416 36576 33468 36582
rect 33416 36518 33468 36524
rect 33152 36378 33180 36518
rect 32128 36372 32180 36378
rect 32128 36314 32180 36320
rect 33140 36372 33192 36378
rect 33140 36314 33192 36320
rect 32140 35698 32168 36314
rect 33428 35834 33456 36518
rect 34520 36168 34572 36174
rect 34520 36110 34572 36116
rect 33416 35828 33468 35834
rect 33416 35770 33468 35776
rect 32128 35692 32180 35698
rect 32128 35634 32180 35640
rect 32588 35692 32640 35698
rect 32588 35634 32640 35640
rect 33692 35692 33744 35698
rect 33692 35634 33744 35640
rect 31392 34944 31444 34950
rect 31392 34886 31444 34892
rect 31116 34740 31168 34746
rect 31116 34682 31168 34688
rect 31128 33862 31156 34682
rect 31404 34610 31432 34886
rect 32140 34678 32168 35634
rect 32600 35290 32628 35634
rect 32588 35284 32640 35290
rect 32588 35226 32640 35232
rect 33232 35080 33284 35086
rect 33232 35022 33284 35028
rect 33244 34746 33272 35022
rect 33232 34740 33284 34746
rect 33232 34682 33284 34688
rect 32128 34672 32180 34678
rect 32128 34614 32180 34620
rect 31392 34604 31444 34610
rect 31392 34546 31444 34552
rect 31760 34400 31812 34406
rect 31760 34342 31812 34348
rect 31772 33998 31800 34342
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31116 33856 31168 33862
rect 31116 33798 31168 33804
rect 31128 33318 31156 33798
rect 31772 33454 31800 33934
rect 32140 33590 32168 34614
rect 33704 34610 33732 35634
rect 33876 35012 33928 35018
rect 33876 34954 33928 34960
rect 33888 34610 33916 34954
rect 34532 34610 34560 36110
rect 34716 35834 34744 37266
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 34808 36258 34836 37198
rect 35256 37188 35308 37194
rect 35452 37176 35480 37402
rect 35532 37324 35584 37330
rect 35532 37266 35584 37272
rect 35308 37148 35480 37176
rect 35256 37130 35308 37136
rect 34888 37120 34940 37126
rect 34888 37062 34940 37068
rect 34900 36854 34928 37062
rect 34888 36848 34940 36854
rect 34888 36790 34940 36796
rect 35348 36780 35400 36786
rect 35348 36722 35400 36728
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34808 36230 34928 36258
rect 34900 35834 34928 36230
rect 34704 35828 34756 35834
rect 34704 35770 34756 35776
rect 34888 35828 34940 35834
rect 34888 35770 34940 35776
rect 35360 35494 35388 36722
rect 34796 35488 34848 35494
rect 34796 35430 34848 35436
rect 35348 35488 35400 35494
rect 35348 35430 35400 35436
rect 33692 34604 33744 34610
rect 33692 34546 33744 34552
rect 33876 34604 33928 34610
rect 33876 34546 33928 34552
rect 34520 34604 34572 34610
rect 34520 34546 34572 34552
rect 33888 34134 33916 34546
rect 34336 34400 34388 34406
rect 34336 34342 34388 34348
rect 33876 34128 33928 34134
rect 33876 34070 33928 34076
rect 33888 33930 33916 34070
rect 34348 33998 34376 34342
rect 34532 34066 34560 34546
rect 34520 34060 34572 34066
rect 34520 34002 34572 34008
rect 34808 33998 34836 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35452 34746 35480 37148
rect 35440 34740 35492 34746
rect 35440 34682 35492 34688
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34336 33992 34388 33998
rect 34336 33934 34388 33940
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 33508 33924 33560 33930
rect 33508 33866 33560 33872
rect 33876 33924 33928 33930
rect 33876 33866 33928 33872
rect 32496 33856 32548 33862
rect 32496 33798 32548 33804
rect 32128 33584 32180 33590
rect 32128 33526 32180 33532
rect 31760 33448 31812 33454
rect 31760 33390 31812 33396
rect 31116 33312 31168 33318
rect 31116 33254 31168 33260
rect 31392 33312 31444 33318
rect 31392 33254 31444 33260
rect 31404 32910 31432 33254
rect 32140 32978 32168 33526
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31760 32836 31812 32842
rect 31760 32778 31812 32784
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 31772 31482 31800 32778
rect 32416 32570 32444 32778
rect 32508 32570 32536 33798
rect 33520 33522 33548 33866
rect 34520 33856 34572 33862
rect 34520 33798 34572 33804
rect 34532 33590 34560 33798
rect 34808 33658 34836 33934
rect 34796 33652 34848 33658
rect 34796 33594 34848 33600
rect 34520 33584 34572 33590
rect 34520 33526 34572 33532
rect 33508 33516 33560 33522
rect 33508 33458 33560 33464
rect 33416 33448 33468 33454
rect 33416 33390 33468 33396
rect 33428 32774 33456 33390
rect 34152 33312 34204 33318
rect 34152 33254 34204 33260
rect 34164 32910 34192 33254
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34152 32904 34204 32910
rect 34152 32846 34204 32852
rect 32772 32768 32824 32774
rect 32772 32710 32824 32716
rect 33416 32768 33468 32774
rect 33416 32710 33468 32716
rect 33968 32768 34020 32774
rect 33968 32710 34020 32716
rect 32404 32564 32456 32570
rect 32404 32506 32456 32512
rect 32496 32564 32548 32570
rect 32496 32506 32548 32512
rect 32784 32502 32812 32710
rect 32772 32496 32824 32502
rect 32772 32438 32824 32444
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32416 31482 32444 32370
rect 32772 32360 32824 32366
rect 32772 32302 32824 32308
rect 31760 31476 31812 31482
rect 31760 31418 31812 31424
rect 32404 31476 32456 31482
rect 32404 31418 32456 31424
rect 32128 31408 32180 31414
rect 32128 31350 32180 31356
rect 32140 31278 32168 31350
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32128 31272 32180 31278
rect 32128 31214 32180 31220
rect 31208 31136 31260 31142
rect 31208 31078 31260 31084
rect 31220 30802 31248 31078
rect 31208 30796 31260 30802
rect 31208 30738 31260 30744
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 31404 30326 31432 30670
rect 31668 30592 31720 30598
rect 31668 30534 31720 30540
rect 31392 30320 31444 30326
rect 31392 30262 31444 30268
rect 31680 30258 31708 30534
rect 32140 30258 32168 31214
rect 32508 31142 32536 31282
rect 32496 31136 32548 31142
rect 32496 31078 32548 31084
rect 32220 30728 32272 30734
rect 32220 30670 32272 30676
rect 31668 30252 31720 30258
rect 31668 30194 31720 30200
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 31576 30048 31628 30054
rect 31576 29990 31628 29996
rect 31588 29646 31616 29990
rect 31576 29640 31628 29646
rect 31576 29582 31628 29588
rect 32232 29510 32260 30670
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 32324 29850 32352 30194
rect 32312 29844 32364 29850
rect 32312 29786 32364 29792
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 32220 29504 32272 29510
rect 32220 29446 32272 29452
rect 30748 29164 30800 29170
rect 30748 29106 30800 29112
rect 30760 28762 30788 29106
rect 30748 28756 30800 28762
rect 30748 28698 30800 28704
rect 31772 28558 31800 29446
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 30656 28484 30708 28490
rect 30656 28426 30708 28432
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 29932 28082 29960 28358
rect 30668 28234 30696 28426
rect 30668 28206 30788 28234
rect 29920 28076 29972 28082
rect 29920 28018 29972 28024
rect 30656 28076 30708 28082
rect 30656 28018 30708 28024
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 29828 27532 29880 27538
rect 29828 27474 29880 27480
rect 29840 26042 29868 27474
rect 30196 27396 30248 27402
rect 30196 27338 30248 27344
rect 30208 27130 30236 27338
rect 30196 27124 30248 27130
rect 30196 27066 30248 27072
rect 30392 27062 30420 27814
rect 30668 27334 30696 28018
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30668 27062 30696 27270
rect 30380 27056 30432 27062
rect 30380 26998 30432 27004
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30668 26858 30696 26998
rect 30656 26852 30708 26858
rect 30656 26794 30708 26800
rect 29828 26036 29880 26042
rect 29828 25978 29880 25984
rect 30760 25838 30788 28206
rect 31024 27124 31076 27130
rect 31024 27066 31076 27072
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 30748 25832 30800 25838
rect 30748 25774 30800 25780
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 29828 25220 29880 25226
rect 29828 25162 29880 25168
rect 29840 24954 29868 25162
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 29828 24948 29880 24954
rect 29828 24890 29880 24896
rect 30392 24750 30420 25094
rect 30748 24880 30800 24886
rect 30748 24822 30800 24828
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 30392 24410 30420 24686
rect 30472 24676 30524 24682
rect 30472 24618 30524 24624
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30484 24206 30512 24618
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 30472 24200 30524 24206
rect 30472 24142 30524 24148
rect 28448 23656 28500 23662
rect 28448 23598 28500 23604
rect 28080 23520 28132 23526
rect 28080 23462 28132 23468
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 27804 23248 27856 23254
rect 27804 23190 27856 23196
rect 27712 23180 27764 23186
rect 27712 23122 27764 23128
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 28172 23112 28224 23118
rect 28172 23054 28224 23060
rect 27816 22982 27844 23054
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27540 22642 27660 22658
rect 27540 22636 27672 22642
rect 27540 22630 27620 22636
rect 27540 22506 27568 22630
rect 27620 22578 27672 22584
rect 27816 22506 27844 22918
rect 28184 22642 28212 23054
rect 28460 22778 28488 23598
rect 28552 23322 28580 24142
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28644 23186 28672 24142
rect 30380 24132 30432 24138
rect 30380 24074 30432 24080
rect 30392 23866 30420 24074
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30380 23860 30432 23866
rect 30380 23802 30432 23808
rect 30484 23730 30512 24006
rect 30564 23860 30616 23866
rect 30564 23802 30616 23808
rect 30472 23724 30524 23730
rect 30472 23666 30524 23672
rect 28632 23180 28684 23186
rect 28632 23122 28684 23128
rect 29920 22976 29972 22982
rect 29920 22918 29972 22924
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 27528 22500 27580 22506
rect 27528 22442 27580 22448
rect 27804 22500 27856 22506
rect 27804 22442 27856 22448
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 26884 21548 26936 21554
rect 26884 21490 26936 21496
rect 26700 20868 26752 20874
rect 26700 20810 26752 20816
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26344 20398 26372 20742
rect 26712 20602 26740 20810
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26988 20398 27016 22170
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 27448 20466 27476 21286
rect 27528 20868 27580 20874
rect 27528 20810 27580 20816
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 26332 20392 26384 20398
rect 26332 20334 26384 20340
rect 26976 20392 27028 20398
rect 26976 20334 27028 20340
rect 27540 20262 27568 20810
rect 28184 20806 28212 22578
rect 29932 22574 29960 22918
rect 30484 22710 30512 23666
rect 30576 23254 30604 23802
rect 30760 23798 30788 24822
rect 30852 24818 30880 25638
rect 30944 25362 30972 25842
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30944 24954 30972 25298
rect 30932 24948 30984 24954
rect 30932 24890 30984 24896
rect 31036 24818 31064 27066
rect 31300 27056 31352 27062
rect 31300 26998 31352 27004
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 31220 25974 31248 26250
rect 31208 25968 31260 25974
rect 31208 25910 31260 25916
rect 31208 25152 31260 25158
rect 31208 25094 31260 25100
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 31024 24812 31076 24818
rect 31024 24754 31076 24760
rect 30748 23792 30800 23798
rect 30748 23734 30800 23740
rect 30932 23792 30984 23798
rect 30932 23734 30984 23740
rect 30564 23248 30616 23254
rect 30616 23196 30788 23202
rect 30564 23190 30788 23196
rect 30576 23174 30788 23190
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30472 22704 30524 22710
rect 30472 22646 30524 22652
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 29920 22568 29972 22574
rect 29920 22510 29972 22516
rect 29460 22432 29512 22438
rect 29460 22374 29512 22380
rect 30392 22386 30420 22578
rect 30668 22506 30696 23054
rect 30760 22710 30788 23174
rect 30944 22930 30972 23734
rect 31220 23662 31248 25094
rect 31312 23866 31340 26998
rect 31772 26586 31800 28494
rect 32312 28416 32364 28422
rect 32312 28358 32364 28364
rect 32324 28082 32352 28358
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 31944 27872 31996 27878
rect 31944 27814 31996 27820
rect 31852 27532 31904 27538
rect 31852 27474 31904 27480
rect 31864 26858 31892 27474
rect 31956 27470 31984 27814
rect 32324 27538 32352 28018
rect 32588 28008 32640 28014
rect 32588 27950 32640 27956
rect 32680 28008 32732 28014
rect 32680 27950 32732 27956
rect 32312 27532 32364 27538
rect 32312 27474 32364 27480
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 31956 27130 31984 27406
rect 31944 27124 31996 27130
rect 31944 27066 31996 27072
rect 31852 26852 31904 26858
rect 31852 26794 31904 26800
rect 31760 26580 31812 26586
rect 31760 26522 31812 26528
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 31588 24410 31616 25230
rect 31772 25226 31800 26522
rect 32600 26246 32628 27950
rect 32692 27606 32720 27950
rect 32680 27600 32732 27606
rect 32680 27542 32732 27548
rect 32588 26240 32640 26246
rect 32588 26182 32640 26188
rect 32496 25696 32548 25702
rect 32496 25638 32548 25644
rect 31760 25220 31812 25226
rect 31760 25162 31812 25168
rect 31772 24818 31800 25162
rect 32508 24886 32536 25638
rect 32600 25362 32628 26182
rect 32588 25356 32640 25362
rect 32588 25298 32640 25304
rect 32496 24880 32548 24886
rect 32496 24822 32548 24828
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31576 24404 31628 24410
rect 31576 24346 31628 24352
rect 31772 24206 31800 24754
rect 31760 24200 31812 24206
rect 31760 24142 31812 24148
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31208 23656 31260 23662
rect 31208 23598 31260 23604
rect 31312 23254 31340 23802
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31300 23248 31352 23254
rect 31300 23190 31352 23196
rect 31300 23112 31352 23118
rect 31300 23054 31352 23060
rect 31116 22976 31168 22982
rect 30944 22924 31116 22930
rect 30944 22918 31168 22924
rect 30944 22902 31156 22918
rect 30748 22704 30800 22710
rect 30748 22646 30800 22652
rect 30944 22642 30972 22902
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 31116 22568 31168 22574
rect 31116 22510 31168 22516
rect 30656 22500 30708 22506
rect 30656 22442 30708 22448
rect 30472 22432 30524 22438
rect 30392 22380 30472 22386
rect 30392 22374 30524 22380
rect 29472 21962 29500 22374
rect 30392 22358 30512 22374
rect 30392 22234 30420 22358
rect 31128 22234 31156 22510
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 31116 22228 31168 22234
rect 31116 22170 31168 22176
rect 30392 22094 30420 22170
rect 30392 22066 30512 22094
rect 29736 22024 29788 22030
rect 29736 21966 29788 21972
rect 29460 21956 29512 21962
rect 29460 21898 29512 21904
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28276 21146 28304 21490
rect 28264 21140 28316 21146
rect 28264 21082 28316 21088
rect 28172 20800 28224 20806
rect 28172 20742 28224 20748
rect 28184 20602 28212 20742
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28276 20466 28304 21082
rect 29748 20942 29776 21966
rect 30196 21684 30248 21690
rect 30196 21626 30248 21632
rect 29920 21344 29972 21350
rect 29920 21286 29972 21292
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29828 20868 29880 20874
rect 29828 20810 29880 20816
rect 29840 20602 29868 20810
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29932 20466 29960 21286
rect 30208 20466 30236 21626
rect 30484 21622 30512 22066
rect 30472 21616 30524 21622
rect 30472 21558 30524 21564
rect 31312 20942 31340 23054
rect 31404 22642 31432 23462
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31484 22636 31536 22642
rect 31484 22578 31536 22584
rect 31404 21690 31432 22578
rect 31392 21684 31444 21690
rect 31392 21626 31444 21632
rect 31404 21146 31432 21626
rect 31496 21554 31524 22578
rect 32508 22438 32536 24822
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31496 21146 31524 21490
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 31484 21140 31536 21146
rect 31484 21082 31536 21088
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31496 20466 31524 21082
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31864 20602 31892 20810
rect 31852 20596 31904 20602
rect 31852 20538 31904 20544
rect 32324 20466 32352 20878
rect 32784 20641 32812 32302
rect 33140 30660 33192 30666
rect 33140 30602 33192 30608
rect 33152 30394 33180 30602
rect 33140 30388 33192 30394
rect 33140 30330 33192 30336
rect 33428 29238 33456 32710
rect 33980 32434 34008 32710
rect 33968 32428 34020 32434
rect 33968 32370 34020 32376
rect 33980 31414 34008 32370
rect 35544 32366 35572 37266
rect 36820 37256 36872 37262
rect 36820 37198 36872 37204
rect 36176 37188 36228 37194
rect 36176 37130 36228 37136
rect 35900 37120 35952 37126
rect 35900 37062 35952 37068
rect 35624 36848 35676 36854
rect 35624 36790 35676 36796
rect 35532 32360 35584 32366
rect 35532 32302 35584 32308
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35636 31890 35664 36790
rect 35912 36106 35940 37062
rect 36188 36922 36216 37130
rect 36452 37120 36504 37126
rect 36452 37062 36504 37068
rect 36176 36916 36228 36922
rect 36176 36858 36228 36864
rect 36464 36786 36492 37062
rect 36728 36848 36780 36854
rect 36728 36790 36780 36796
rect 36452 36780 36504 36786
rect 36452 36722 36504 36728
rect 35900 36100 35952 36106
rect 35900 36042 35952 36048
rect 35912 35834 35940 36042
rect 36740 36038 36768 36790
rect 36832 36038 36860 37198
rect 36728 36032 36780 36038
rect 36728 35974 36780 35980
rect 36820 36032 36872 36038
rect 36820 35974 36872 35980
rect 35900 35828 35952 35834
rect 35900 35770 35952 35776
rect 35716 34604 35768 34610
rect 35716 34546 35768 34552
rect 35728 34202 35756 34546
rect 35716 34196 35768 34202
rect 35716 34138 35768 34144
rect 36740 32026 36768 35974
rect 36832 35766 36860 35974
rect 36820 35760 36872 35766
rect 36820 35702 36872 35708
rect 37108 34406 37136 38286
rect 37200 37262 37228 38354
rect 37464 37800 37516 37806
rect 37464 37742 37516 37748
rect 37476 37670 37504 37742
rect 37464 37664 37516 37670
rect 37464 37606 37516 37612
rect 37280 37460 37332 37466
rect 37280 37402 37332 37408
rect 37188 37256 37240 37262
rect 37188 37198 37240 37204
rect 37200 36242 37228 37198
rect 37292 36718 37320 37402
rect 37476 36922 37504 37606
rect 37568 37194 37596 38898
rect 38120 37670 38148 39374
rect 38660 39296 38712 39302
rect 38660 39238 38712 39244
rect 38108 37664 38160 37670
rect 38108 37606 38160 37612
rect 37924 37460 37976 37466
rect 37924 37402 37976 37408
rect 37556 37188 37608 37194
rect 37556 37130 37608 37136
rect 37464 36916 37516 36922
rect 37464 36858 37516 36864
rect 37280 36712 37332 36718
rect 37280 36654 37332 36660
rect 37188 36236 37240 36242
rect 37188 36178 37240 36184
rect 37476 36174 37504 36858
rect 37568 36786 37596 37130
rect 37556 36780 37608 36786
rect 37556 36722 37608 36728
rect 37464 36168 37516 36174
rect 37464 36110 37516 36116
rect 37096 34400 37148 34406
rect 37096 34342 37148 34348
rect 37108 33590 37136 34342
rect 37464 33924 37516 33930
rect 37464 33866 37516 33872
rect 37476 33658 37504 33866
rect 37464 33652 37516 33658
rect 37464 33594 37516 33600
rect 37096 33584 37148 33590
rect 37096 33526 37148 33532
rect 36728 32020 36780 32026
rect 36728 31962 36780 31968
rect 37108 31958 37136 33526
rect 37568 33522 37596 36722
rect 37832 36576 37884 36582
rect 37832 36518 37884 36524
rect 37844 35698 37872 36518
rect 37832 35692 37884 35698
rect 37832 35634 37884 35640
rect 37740 34060 37792 34066
rect 37740 34002 37792 34008
rect 37752 33522 37780 34002
rect 37556 33516 37608 33522
rect 37556 33458 37608 33464
rect 37740 33516 37792 33522
rect 37740 33458 37792 33464
rect 37188 32836 37240 32842
rect 37188 32778 37240 32784
rect 37280 32836 37332 32842
rect 37280 32778 37332 32784
rect 37200 32298 37228 32778
rect 37188 32292 37240 32298
rect 37188 32234 37240 32240
rect 37188 32020 37240 32026
rect 37188 31962 37240 31968
rect 37096 31952 37148 31958
rect 37096 31894 37148 31900
rect 35624 31884 35676 31890
rect 35624 31826 35676 31832
rect 33968 31408 34020 31414
rect 33968 31350 34020 31356
rect 34060 31272 34112 31278
rect 34060 31214 34112 31220
rect 33600 31204 33652 31210
rect 33600 31146 33652 31152
rect 33612 30938 33640 31146
rect 33600 30932 33652 30938
rect 33600 30874 33652 30880
rect 34072 30734 34100 31214
rect 35440 31136 35492 31142
rect 35440 31078 35492 31084
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34060 30728 34112 30734
rect 34060 30670 34112 30676
rect 35452 30258 35480 31078
rect 35440 30252 35492 30258
rect 35440 30194 35492 30200
rect 35348 30048 35400 30054
rect 35348 29990 35400 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34244 29640 34296 29646
rect 34244 29582 34296 29588
rect 34256 29238 34284 29582
rect 34612 29572 34664 29578
rect 34612 29514 34664 29520
rect 33416 29232 33468 29238
rect 33416 29174 33468 29180
rect 34244 29232 34296 29238
rect 34244 29174 34296 29180
rect 34624 29034 34652 29514
rect 35360 29170 35388 29990
rect 35452 29782 35480 30194
rect 35440 29776 35492 29782
rect 35440 29718 35492 29724
rect 35636 29578 35664 31826
rect 35900 31816 35952 31822
rect 35900 31758 35952 31764
rect 36084 31816 36136 31822
rect 36084 31758 36136 31764
rect 35912 31346 35940 31758
rect 35900 31340 35952 31346
rect 35900 31282 35952 31288
rect 35900 31136 35952 31142
rect 35900 31078 35952 31084
rect 35912 30666 35940 31078
rect 35900 30660 35952 30666
rect 35900 30602 35952 30608
rect 35624 29572 35676 29578
rect 35676 29532 35756 29560
rect 35624 29514 35676 29520
rect 35728 29306 35756 29532
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 35716 29300 35768 29306
rect 35716 29242 35768 29248
rect 35348 29164 35400 29170
rect 35400 29124 35664 29152
rect 35348 29106 35400 29112
rect 34612 29028 34664 29034
rect 34612 28970 34664 28976
rect 34704 28960 34756 28966
rect 34704 28902 34756 28908
rect 35256 28960 35308 28966
rect 35308 28908 35388 28914
rect 35256 28902 35388 28908
rect 34716 28490 34744 28902
rect 35268 28886 35388 28902
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 32956 28484 33008 28490
rect 32956 28426 33008 28432
rect 34704 28484 34756 28490
rect 34704 28426 34756 28432
rect 32968 28218 32996 28426
rect 32956 28212 33008 28218
rect 32956 28154 33008 28160
rect 34796 27872 34848 27878
rect 34796 27814 34848 27820
rect 33784 27600 33836 27606
rect 33784 27542 33836 27548
rect 33692 27396 33744 27402
rect 33692 27338 33744 27344
rect 33704 26994 33732 27338
rect 33796 27334 33824 27542
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 33508 26988 33560 26994
rect 33508 26930 33560 26936
rect 33692 26988 33744 26994
rect 33692 26930 33744 26936
rect 32956 26920 33008 26926
rect 32956 26862 33008 26868
rect 32968 26586 32996 26862
rect 33520 26586 33548 26930
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 33508 26580 33560 26586
rect 33508 26522 33560 26528
rect 33704 25974 33732 26930
rect 33692 25968 33744 25974
rect 33692 25910 33744 25916
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 32968 24274 32996 24754
rect 33796 24698 33824 27270
rect 34808 26976 34836 27814
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27470 35388 28886
rect 35440 28620 35492 28626
rect 35440 28562 35492 28568
rect 35452 28014 35480 28562
rect 35636 28558 35664 29124
rect 35912 29102 35940 29446
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 35900 29096 35952 29102
rect 35900 29038 35952 29044
rect 35912 28558 35940 29038
rect 36004 28762 36032 29106
rect 35992 28756 36044 28762
rect 35992 28698 36044 28704
rect 35992 28620 36044 28626
rect 35992 28562 36044 28568
rect 35624 28552 35676 28558
rect 35624 28494 35676 28500
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35532 28416 35584 28422
rect 35532 28358 35584 28364
rect 35440 28008 35492 28014
rect 35440 27950 35492 27956
rect 35544 27538 35572 28358
rect 35636 27946 35664 28494
rect 36004 28082 36032 28562
rect 35992 28076 36044 28082
rect 35992 28018 36044 28024
rect 35624 27940 35676 27946
rect 35624 27882 35676 27888
rect 35532 27532 35584 27538
rect 35532 27474 35584 27480
rect 35348 27464 35400 27470
rect 35348 27406 35400 27412
rect 35348 27328 35400 27334
rect 35348 27270 35400 27276
rect 35360 27130 35388 27270
rect 35348 27124 35400 27130
rect 35348 27066 35400 27072
rect 35072 26988 35124 26994
rect 34808 26948 35072 26976
rect 35072 26930 35124 26936
rect 35084 26790 35112 26930
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 35072 26784 35124 26790
rect 35072 26726 35124 26732
rect 34808 26450 34836 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34796 26444 34848 26450
rect 34796 26386 34848 26392
rect 35360 26382 35388 27066
rect 35440 26444 35492 26450
rect 35440 26386 35492 26392
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 25362 35388 26318
rect 35452 26042 35480 26386
rect 35440 26036 35492 26042
rect 35440 25978 35492 25984
rect 35544 25906 35572 27474
rect 35900 27396 35952 27402
rect 35900 27338 35952 27344
rect 35532 25900 35584 25906
rect 35532 25842 35584 25848
rect 35348 25356 35400 25362
rect 35348 25298 35400 25304
rect 35624 25220 35676 25226
rect 35624 25162 35676 25168
rect 34796 24880 34848 24886
rect 34796 24822 34848 24828
rect 33704 24670 33824 24698
rect 32956 24268 33008 24274
rect 32956 24210 33008 24216
rect 32968 22624 32996 24210
rect 33704 23730 33732 24670
rect 34808 24206 34836 24822
rect 35440 24812 35492 24818
rect 35440 24754 35492 24760
rect 35348 24608 35400 24614
rect 35348 24550 35400 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24206 35388 24550
rect 35452 24410 35480 24754
rect 35440 24404 35492 24410
rect 35440 24346 35492 24352
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 35348 24200 35400 24206
rect 35348 24142 35400 24148
rect 33784 24132 33836 24138
rect 33784 24074 33836 24080
rect 33796 23866 33824 24074
rect 34612 24064 34664 24070
rect 34612 24006 34664 24012
rect 33784 23860 33836 23866
rect 33784 23802 33836 23808
rect 34624 23730 34652 24006
rect 35360 23798 35388 24142
rect 35348 23792 35400 23798
rect 35348 23734 35400 23740
rect 33692 23724 33744 23730
rect 33692 23666 33744 23672
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 33704 23118 33732 23666
rect 33692 23112 33744 23118
rect 33692 23054 33744 23060
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 33140 22636 33192 22642
rect 32968 22596 33140 22624
rect 33060 20942 33088 22596
rect 33140 22578 33192 22584
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33888 22234 33916 22578
rect 33876 22228 33928 22234
rect 33876 22170 33928 22176
rect 33980 21962 34008 23054
rect 34624 23050 34652 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34704 23316 34756 23322
rect 34704 23258 34756 23264
rect 34612 23044 34664 23050
rect 34612 22986 34664 22992
rect 34624 21962 34652 22986
rect 34716 22438 34744 23258
rect 34796 23248 34848 23254
rect 34796 23190 34848 23196
rect 34704 22432 34756 22438
rect 34704 22374 34756 22380
rect 34716 22030 34744 22374
rect 34808 22098 34836 23190
rect 35360 23050 35388 23734
rect 35348 23044 35400 23050
rect 35348 22986 35400 22992
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22092 34848 22098
rect 34796 22034 34848 22040
rect 35360 22030 35388 22986
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 33968 21956 34020 21962
rect 33968 21898 34020 21904
rect 34336 21956 34388 21962
rect 34336 21898 34388 21904
rect 34612 21956 34664 21962
rect 34612 21898 34664 21904
rect 33048 20936 33100 20942
rect 33048 20878 33100 20884
rect 32770 20632 32826 20641
rect 32770 20567 32826 20576
rect 34348 20534 34376 21898
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 34610 20632 34666 20641
rect 35360 20602 35388 20810
rect 34610 20567 34666 20576
rect 35348 20596 35400 20602
rect 34336 20528 34388 20534
rect 34336 20470 34388 20476
rect 34624 20466 34652 20567
rect 35348 20538 35400 20544
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 31484 20460 31536 20466
rect 31484 20402 31536 20408
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 34612 20460 34664 20466
rect 34612 20402 34664 20408
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 32876 20058 32904 20402
rect 33506 20360 33562 20369
rect 33506 20295 33562 20304
rect 33048 20256 33100 20262
rect 33048 20198 33100 20204
rect 32864 20052 32916 20058
rect 32864 19994 32916 20000
rect 33060 19378 33088 20198
rect 33324 19848 33376 19854
rect 33324 19790 33376 19796
rect 33336 19514 33364 19790
rect 33324 19508 33376 19514
rect 33324 19450 33376 19456
rect 33048 19372 33100 19378
rect 33048 19314 33100 19320
rect 33520 19310 33548 20295
rect 33692 20256 33744 20262
rect 33692 20198 33744 20204
rect 33704 19922 33732 20198
rect 33692 19916 33744 19922
rect 33692 19858 33744 19864
rect 33888 19786 33916 20402
rect 34244 20256 34296 20262
rect 34244 20198 34296 20204
rect 33968 20052 34020 20058
rect 33968 19994 34020 20000
rect 33980 19961 34008 19994
rect 34256 19990 34284 20198
rect 34808 20058 34836 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34796 20052 34848 20058
rect 34796 19994 34848 20000
rect 34244 19984 34296 19990
rect 33966 19952 34022 19961
rect 34244 19926 34296 19932
rect 35346 19952 35402 19961
rect 33966 19887 34022 19896
rect 33876 19780 33928 19786
rect 33876 19722 33928 19728
rect 33980 19310 34008 19887
rect 33508 19304 33560 19310
rect 33508 19246 33560 19252
rect 33968 19304 34020 19310
rect 33968 19246 34020 19252
rect 34256 18766 34284 19926
rect 35346 19887 35402 19896
rect 35360 19854 35388 19887
rect 34612 19848 34664 19854
rect 34610 19816 34612 19825
rect 35348 19848 35400 19854
rect 34664 19816 34666 19825
rect 34336 19780 34388 19786
rect 34716 19786 34928 19802
rect 35348 19790 35400 19796
rect 34610 19751 34666 19760
rect 34704 19780 34928 19786
rect 34336 19722 34388 19728
rect 34756 19774 34928 19780
rect 34704 19722 34756 19728
rect 34348 18970 34376 19722
rect 34796 19712 34848 19718
rect 34900 19700 34928 19774
rect 34980 19712 35032 19718
rect 34900 19672 34980 19700
rect 34796 19654 34848 19660
rect 34980 19654 35032 19660
rect 34808 19428 34836 19654
rect 35164 19508 35216 19514
rect 35164 19450 35216 19456
rect 35440 19508 35492 19514
rect 35440 19450 35492 19456
rect 34980 19440 35032 19446
rect 34808 19400 34980 19428
rect 34980 19382 35032 19388
rect 35176 19310 35204 19450
rect 35164 19304 35216 19310
rect 35164 19246 35216 19252
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 34244 18760 34296 18766
rect 34244 18702 34296 18708
rect 35452 18426 35480 19450
rect 35636 18834 35664 25162
rect 35716 24744 35768 24750
rect 35716 24686 35768 24692
rect 35728 24410 35756 24686
rect 35716 24404 35768 24410
rect 35716 24346 35768 24352
rect 35728 24070 35756 24346
rect 35716 24064 35768 24070
rect 35716 24006 35768 24012
rect 35912 22094 35940 27338
rect 36096 24614 36124 31758
rect 36176 30592 36228 30598
rect 36176 30534 36228 30540
rect 36188 30326 36216 30534
rect 36176 30320 36228 30326
rect 36176 30262 36228 30268
rect 36188 29646 36216 30262
rect 36176 29640 36228 29646
rect 36176 29582 36228 29588
rect 36360 29504 36412 29510
rect 36360 29446 36412 29452
rect 36372 28694 36400 29446
rect 36636 28960 36688 28966
rect 36636 28902 36688 28908
rect 36360 28688 36412 28694
rect 36360 28630 36412 28636
rect 36268 28416 36320 28422
rect 36268 28358 36320 28364
rect 36176 26988 36228 26994
rect 36176 26930 36228 26936
rect 36188 26042 36216 26930
rect 36176 26036 36228 26042
rect 36176 25978 36228 25984
rect 36176 25288 36228 25294
rect 36176 25230 36228 25236
rect 36084 24608 36136 24614
rect 36084 24550 36136 24556
rect 35992 24132 36044 24138
rect 35992 24074 36044 24080
rect 36004 23730 36032 24074
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 35912 22066 36032 22094
rect 35808 20460 35860 20466
rect 35808 20402 35860 20408
rect 35820 20058 35848 20402
rect 36004 20262 36032 22066
rect 36084 20460 36136 20466
rect 36084 20402 36136 20408
rect 36096 20369 36124 20402
rect 36082 20360 36138 20369
rect 36082 20295 36138 20304
rect 35992 20256 36044 20262
rect 35992 20198 36044 20204
rect 35808 20052 35860 20058
rect 35808 19994 35860 20000
rect 35900 20052 35952 20058
rect 35900 19994 35952 20000
rect 35912 19854 35940 19994
rect 35900 19848 35952 19854
rect 35900 19790 35952 19796
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35716 19440 35768 19446
rect 35716 19382 35768 19388
rect 35728 18970 35756 19382
rect 35820 19378 35848 19654
rect 36004 19446 36032 20198
rect 36188 20058 36216 25230
rect 36280 25226 36308 28358
rect 36372 28150 36400 28630
rect 36648 28558 36676 28902
rect 36912 28756 36964 28762
rect 36912 28698 36964 28704
rect 36636 28552 36688 28558
rect 36636 28494 36688 28500
rect 36360 28144 36412 28150
rect 36360 28086 36412 28092
rect 36924 27130 36952 28698
rect 36912 27124 36964 27130
rect 36912 27066 36964 27072
rect 36728 26852 36780 26858
rect 36728 26794 36780 26800
rect 36544 26580 36596 26586
rect 36544 26522 36596 26528
rect 36556 26042 36584 26522
rect 36740 26314 36768 26794
rect 36728 26308 36780 26314
rect 36728 26250 36780 26256
rect 36820 26308 36872 26314
rect 36820 26250 36872 26256
rect 36544 26036 36596 26042
rect 36544 25978 36596 25984
rect 36360 25900 36412 25906
rect 36360 25842 36412 25848
rect 36728 25900 36780 25906
rect 36832 25888 36860 26250
rect 36780 25860 36860 25888
rect 36728 25842 36780 25848
rect 36372 25498 36400 25842
rect 36360 25492 36412 25498
rect 36360 25434 36412 25440
rect 36268 25220 36320 25226
rect 36268 25162 36320 25168
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36280 22574 36308 23666
rect 36372 22642 36400 23666
rect 36636 23520 36688 23526
rect 36636 23462 36688 23468
rect 36648 23118 36676 23462
rect 36636 23112 36688 23118
rect 36636 23054 36688 23060
rect 36636 22704 36688 22710
rect 36636 22646 36688 22652
rect 36360 22636 36412 22642
rect 36360 22578 36412 22584
rect 36544 22636 36596 22642
rect 36544 22578 36596 22584
rect 36268 22568 36320 22574
rect 36268 22510 36320 22516
rect 36268 20800 36320 20806
rect 36268 20742 36320 20748
rect 36280 20398 36308 20742
rect 36360 20460 36412 20466
rect 36360 20402 36412 20408
rect 36268 20392 36320 20398
rect 36268 20334 36320 20340
rect 36176 20052 36228 20058
rect 36176 19994 36228 20000
rect 35992 19440 36044 19446
rect 35992 19382 36044 19388
rect 35808 19372 35860 19378
rect 35808 19314 35860 19320
rect 35716 18964 35768 18970
rect 35716 18906 35768 18912
rect 36188 18834 36216 19994
rect 36280 19922 36308 20334
rect 36268 19916 36320 19922
rect 36268 19858 36320 19864
rect 36372 19514 36400 20402
rect 36556 20262 36584 22578
rect 36648 22234 36676 22646
rect 36636 22228 36688 22234
rect 36636 22170 36688 22176
rect 36544 20256 36596 20262
rect 36544 20198 36596 20204
rect 36360 19508 36412 19514
rect 36360 19450 36412 19456
rect 35624 18828 35676 18834
rect 35624 18770 35676 18776
rect 36176 18828 36228 18834
rect 36176 18770 36228 18776
rect 35440 18420 35492 18426
rect 35440 18362 35492 18368
rect 35636 18222 35664 18770
rect 36556 18766 36584 20198
rect 36740 19825 36768 25842
rect 36924 25838 36952 27066
rect 37200 26858 37228 31962
rect 37292 30716 37320 32778
rect 37740 32768 37792 32774
rect 37740 32710 37792 32716
rect 37464 32428 37516 32434
rect 37464 32370 37516 32376
rect 37556 32428 37608 32434
rect 37556 32370 37608 32376
rect 37476 32026 37504 32370
rect 37464 32020 37516 32026
rect 37464 31962 37516 31968
rect 37464 31884 37516 31890
rect 37464 31826 37516 31832
rect 37476 31346 37504 31826
rect 37568 31482 37596 32370
rect 37752 31890 37780 32710
rect 37740 31884 37792 31890
rect 37740 31826 37792 31832
rect 37556 31476 37608 31482
rect 37556 31418 37608 31424
rect 37464 31340 37516 31346
rect 37464 31282 37516 31288
rect 37464 30728 37516 30734
rect 37292 30688 37464 30716
rect 37464 30670 37516 30676
rect 37476 29102 37504 30670
rect 37464 29096 37516 29102
rect 37464 29038 37516 29044
rect 37188 26852 37240 26858
rect 37188 26794 37240 26800
rect 37832 26784 37884 26790
rect 37832 26726 37884 26732
rect 37188 26512 37240 26518
rect 37188 26454 37240 26460
rect 37200 25906 37228 26454
rect 37844 25906 37872 26726
rect 37936 26246 37964 37402
rect 38672 37346 38700 39238
rect 38764 38350 38792 42094
rect 40224 42016 40276 42022
rect 40224 41958 40276 41964
rect 40236 41138 40264 41958
rect 40224 41132 40276 41138
rect 40224 41074 40276 41080
rect 41788 41132 41840 41138
rect 41788 41074 41840 41080
rect 39580 40996 39632 41002
rect 39580 40938 39632 40944
rect 39592 40526 39620 40938
rect 39672 40928 39724 40934
rect 39672 40870 39724 40876
rect 41144 40928 41196 40934
rect 41144 40870 41196 40876
rect 39580 40520 39632 40526
rect 39580 40462 39632 40468
rect 39212 40384 39264 40390
rect 39212 40326 39264 40332
rect 39224 40118 39252 40326
rect 39212 40112 39264 40118
rect 39212 40054 39264 40060
rect 39684 39438 39712 40870
rect 41156 40526 41184 40870
rect 40224 40520 40276 40526
rect 40224 40462 40276 40468
rect 41144 40520 41196 40526
rect 41144 40462 41196 40468
rect 39672 39432 39724 39438
rect 39672 39374 39724 39380
rect 40236 39098 40264 40462
rect 41604 40452 41656 40458
rect 41604 40394 41656 40400
rect 41616 40050 41644 40394
rect 41800 40050 41828 41074
rect 42248 41064 42300 41070
rect 42248 41006 42300 41012
rect 42260 40730 42288 41006
rect 42524 40928 42576 40934
rect 42524 40870 42576 40876
rect 42248 40724 42300 40730
rect 42248 40666 42300 40672
rect 42260 40118 42288 40666
rect 42248 40112 42300 40118
rect 42248 40054 42300 40060
rect 41604 40044 41656 40050
rect 41604 39986 41656 39992
rect 41788 40044 41840 40050
rect 41788 39986 41840 39992
rect 42536 39438 42564 40870
rect 42628 40526 42656 42094
rect 43456 41818 43484 42162
rect 43996 42016 44048 42022
rect 43996 41958 44048 41964
rect 43444 41812 43496 41818
rect 43444 41754 43496 41760
rect 43168 41676 43220 41682
rect 43168 41618 43220 41624
rect 42892 41608 42944 41614
rect 42892 41550 42944 41556
rect 42904 41206 42932 41550
rect 42892 41200 42944 41206
rect 42812 41148 42892 41154
rect 42812 41142 42944 41148
rect 42812 41126 42932 41142
rect 43076 41132 43128 41138
rect 42616 40520 42668 40526
rect 42616 40462 42668 40468
rect 42812 40458 42840 41126
rect 43076 41074 43128 41080
rect 42892 41064 42944 41070
rect 42892 41006 42944 41012
rect 42800 40452 42852 40458
rect 42800 40394 42852 40400
rect 42904 40390 42932 41006
rect 42984 40452 43036 40458
rect 42984 40394 43036 40400
rect 42892 40384 42944 40390
rect 42892 40326 42944 40332
rect 42904 40186 42932 40326
rect 42892 40180 42944 40186
rect 42892 40122 42944 40128
rect 42800 39840 42852 39846
rect 42800 39782 42852 39788
rect 42524 39432 42576 39438
rect 42524 39374 42576 39380
rect 40224 39092 40276 39098
rect 40224 39034 40276 39040
rect 39028 38956 39080 38962
rect 39028 38898 39080 38904
rect 39040 38350 39068 38898
rect 40040 38548 40092 38554
rect 40040 38490 40092 38496
rect 38752 38344 38804 38350
rect 38752 38286 38804 38292
rect 39028 38344 39080 38350
rect 39028 38286 39080 38292
rect 39948 38208 40000 38214
rect 39948 38150 40000 38156
rect 38580 37318 38700 37346
rect 38580 36718 38608 37318
rect 39960 37194 39988 38150
rect 40052 37942 40080 38490
rect 42812 38350 42840 39782
rect 42996 39642 43024 40394
rect 43088 39982 43116 41074
rect 43180 41002 43208 41618
rect 44008 41138 44036 41958
rect 45560 41608 45612 41614
rect 45560 41550 45612 41556
rect 44088 41540 44140 41546
rect 44088 41482 44140 41488
rect 43996 41132 44048 41138
rect 43996 41074 44048 41080
rect 43168 40996 43220 41002
rect 43168 40938 43220 40944
rect 43180 40118 43208 40938
rect 43260 40928 43312 40934
rect 43260 40870 43312 40876
rect 43168 40112 43220 40118
rect 43168 40054 43220 40060
rect 43076 39976 43128 39982
rect 43076 39918 43128 39924
rect 42984 39636 43036 39642
rect 42984 39578 43036 39584
rect 43272 39030 43300 40870
rect 44100 40594 44128 41482
rect 45192 41472 45244 41478
rect 45192 41414 45244 41420
rect 45204 41206 45232 41414
rect 45192 41200 45244 41206
rect 45192 41142 45244 41148
rect 44732 41132 44784 41138
rect 44732 41074 44784 41080
rect 44088 40588 44140 40594
rect 44088 40530 44140 40536
rect 44100 40050 44128 40530
rect 44744 40526 44772 41074
rect 45572 40730 45600 41550
rect 45560 40724 45612 40730
rect 45560 40666 45612 40672
rect 44732 40520 44784 40526
rect 44732 40462 44784 40468
rect 45284 40520 45336 40526
rect 45284 40462 45336 40468
rect 44088 40044 44140 40050
rect 44088 39986 44140 39992
rect 43260 39024 43312 39030
rect 43260 38966 43312 38972
rect 43536 38888 43588 38894
rect 43536 38830 43588 38836
rect 43076 38412 43128 38418
rect 43076 38354 43128 38360
rect 43352 38412 43404 38418
rect 43352 38354 43404 38360
rect 42800 38344 42852 38350
rect 42800 38286 42852 38292
rect 42892 38276 42944 38282
rect 42892 38218 42944 38224
rect 40040 37936 40092 37942
rect 40040 37878 40092 37884
rect 42904 37670 42932 38218
rect 43088 37806 43116 38354
rect 43364 37806 43392 38354
rect 43076 37800 43128 37806
rect 43076 37742 43128 37748
rect 43352 37800 43404 37806
rect 43352 37742 43404 37748
rect 40316 37664 40368 37670
rect 40316 37606 40368 37612
rect 41052 37664 41104 37670
rect 41052 37606 41104 37612
rect 42892 37664 42944 37670
rect 42892 37606 42944 37612
rect 40328 37262 40356 37606
rect 41064 37330 41092 37606
rect 42904 37482 42932 37606
rect 42812 37466 42932 37482
rect 42800 37460 42932 37466
rect 42852 37454 42932 37460
rect 42800 37402 42852 37408
rect 41052 37324 41104 37330
rect 41052 37266 41104 37272
rect 40040 37256 40092 37262
rect 40040 37198 40092 37204
rect 40316 37256 40368 37262
rect 40316 37198 40368 37204
rect 39948 37188 40000 37194
rect 39948 37130 40000 37136
rect 39028 36848 39080 36854
rect 39028 36790 39080 36796
rect 39212 36848 39264 36854
rect 39212 36790 39264 36796
rect 38568 36712 38620 36718
rect 38568 36654 38620 36660
rect 39040 36242 39068 36790
rect 39224 36378 39252 36790
rect 39672 36576 39724 36582
rect 39672 36518 39724 36524
rect 39212 36372 39264 36378
rect 39212 36314 39264 36320
rect 39028 36236 39080 36242
rect 39028 36178 39080 36184
rect 39580 36032 39632 36038
rect 39580 35974 39632 35980
rect 39488 35828 39540 35834
rect 39488 35770 39540 35776
rect 39500 35698 39528 35770
rect 39592 35698 39620 35974
rect 39304 35692 39356 35698
rect 39304 35634 39356 35640
rect 39488 35692 39540 35698
rect 39488 35634 39540 35640
rect 39580 35692 39632 35698
rect 39580 35634 39632 35640
rect 39316 35494 39344 35634
rect 39684 35630 39712 36518
rect 39960 36310 39988 37130
rect 40052 36310 40080 37198
rect 40328 36718 40356 37198
rect 40960 37120 41012 37126
rect 40960 37062 41012 37068
rect 40316 36712 40368 36718
rect 40316 36654 40368 36660
rect 39948 36304 40000 36310
rect 39948 36246 40000 36252
rect 40040 36304 40092 36310
rect 40040 36246 40092 36252
rect 39960 36174 39988 36246
rect 39948 36168 40000 36174
rect 39948 36110 40000 36116
rect 40500 36032 40552 36038
rect 40500 35974 40552 35980
rect 40684 36032 40736 36038
rect 40684 35974 40736 35980
rect 40512 35766 40540 35974
rect 40696 35834 40724 35974
rect 40684 35828 40736 35834
rect 40684 35770 40736 35776
rect 40500 35760 40552 35766
rect 40500 35702 40552 35708
rect 39672 35624 39724 35630
rect 40512 35578 40540 35702
rect 40696 35698 40724 35770
rect 40972 35698 41000 37062
rect 41064 36786 41092 37266
rect 43364 37262 43392 37742
rect 43352 37256 43404 37262
rect 43352 37198 43404 37204
rect 41420 37188 41472 37194
rect 41420 37130 41472 37136
rect 42616 37188 42668 37194
rect 42616 37130 42668 37136
rect 41052 36780 41104 36786
rect 41052 36722 41104 36728
rect 41064 36174 41092 36722
rect 41144 36712 41196 36718
rect 41144 36654 41196 36660
rect 41156 36174 41184 36654
rect 41052 36168 41104 36174
rect 41052 36110 41104 36116
rect 41144 36168 41196 36174
rect 41144 36110 41196 36116
rect 41328 35828 41380 35834
rect 41328 35770 41380 35776
rect 40684 35692 40736 35698
rect 40684 35634 40736 35640
rect 40960 35692 41012 35698
rect 40960 35634 41012 35640
rect 41052 35692 41104 35698
rect 41052 35634 41104 35640
rect 39672 35566 39724 35572
rect 40420 35550 40540 35578
rect 38568 35488 38620 35494
rect 38568 35430 38620 35436
rect 39304 35488 39356 35494
rect 39304 35430 39356 35436
rect 40040 35488 40092 35494
rect 40040 35430 40092 35436
rect 38580 35086 38608 35430
rect 38568 35080 38620 35086
rect 38568 35022 38620 35028
rect 39120 35012 39172 35018
rect 39120 34954 39172 34960
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 38028 34474 38056 34886
rect 38292 34604 38344 34610
rect 38292 34546 38344 34552
rect 38752 34604 38804 34610
rect 38752 34546 38804 34552
rect 38016 34468 38068 34474
rect 38016 34410 38068 34416
rect 38028 33658 38056 34410
rect 38304 34134 38332 34546
rect 38292 34128 38344 34134
rect 38292 34070 38344 34076
rect 38200 33856 38252 33862
rect 38200 33798 38252 33804
rect 38016 33652 38068 33658
rect 38016 33594 38068 33600
rect 38212 33590 38240 33798
rect 38200 33584 38252 33590
rect 38200 33526 38252 33532
rect 38304 33522 38332 34070
rect 38764 33522 38792 34546
rect 38936 34536 38988 34542
rect 38936 34478 38988 34484
rect 38844 34468 38896 34474
rect 38844 34410 38896 34416
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 38752 33516 38804 33522
rect 38752 33458 38804 33464
rect 38660 32768 38712 32774
rect 38660 32710 38712 32716
rect 38384 31816 38436 31822
rect 38304 31764 38384 31770
rect 38304 31758 38436 31764
rect 38304 31742 38424 31758
rect 38568 31748 38620 31754
rect 38108 31136 38160 31142
rect 38108 31078 38160 31084
rect 38120 30734 38148 31078
rect 38108 30728 38160 30734
rect 38108 30670 38160 30676
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 38028 28218 38056 29106
rect 38016 28212 38068 28218
rect 38016 28154 38068 28160
rect 38016 28076 38068 28082
rect 38016 28018 38068 28024
rect 38028 27606 38056 28018
rect 38016 27600 38068 27606
rect 38016 27542 38068 27548
rect 38304 27062 38332 31742
rect 38568 31690 38620 31696
rect 38580 31210 38608 31690
rect 38672 31346 38700 32710
rect 38764 31958 38792 33458
rect 38752 31952 38804 31958
rect 38752 31894 38804 31900
rect 38856 31822 38884 34410
rect 38948 33998 38976 34478
rect 38936 33992 38988 33998
rect 38936 33934 38988 33940
rect 39028 33992 39080 33998
rect 39028 33934 39080 33940
rect 39040 33658 39068 33934
rect 39132 33930 39160 34954
rect 40052 34678 40080 35430
rect 40420 35086 40448 35550
rect 40500 35488 40552 35494
rect 40500 35430 40552 35436
rect 40408 35080 40460 35086
rect 40408 35022 40460 35028
rect 40132 34944 40184 34950
rect 40132 34886 40184 34892
rect 40144 34678 40172 34886
rect 40040 34672 40092 34678
rect 40040 34614 40092 34620
rect 40132 34672 40184 34678
rect 40132 34614 40184 34620
rect 39396 34536 39448 34542
rect 39396 34478 39448 34484
rect 39120 33924 39172 33930
rect 39120 33866 39172 33872
rect 39028 33652 39080 33658
rect 39028 33594 39080 33600
rect 38936 33448 38988 33454
rect 38936 33390 38988 33396
rect 38844 31816 38896 31822
rect 38844 31758 38896 31764
rect 38844 31476 38896 31482
rect 38844 31418 38896 31424
rect 38660 31340 38712 31346
rect 38660 31282 38712 31288
rect 38752 31340 38804 31346
rect 38752 31282 38804 31288
rect 38568 31204 38620 31210
rect 38568 31146 38620 31152
rect 38764 29238 38792 31282
rect 38856 30258 38884 31418
rect 38948 31346 38976 33390
rect 39132 33114 39160 33866
rect 39120 33108 39172 33114
rect 39120 33050 39172 33056
rect 39132 32502 39160 33050
rect 39120 32496 39172 32502
rect 39120 32438 39172 32444
rect 39212 32428 39264 32434
rect 39212 32370 39264 32376
rect 39224 31686 39252 32370
rect 39408 31822 39436 34478
rect 40052 33998 40080 34614
rect 40040 33992 40092 33998
rect 40040 33934 40092 33940
rect 40144 33810 40172 34614
rect 40512 34610 40540 35430
rect 40696 35086 40724 35634
rect 40972 35154 41000 35634
rect 41064 35562 41092 35634
rect 41052 35556 41104 35562
rect 41052 35498 41104 35504
rect 40960 35148 41012 35154
rect 40960 35090 41012 35096
rect 40684 35080 40736 35086
rect 40684 35022 40736 35028
rect 40500 34604 40552 34610
rect 40500 34546 40552 34552
rect 40684 34400 40736 34406
rect 40684 34342 40736 34348
rect 40696 33998 40724 34342
rect 41064 33998 41092 35498
rect 41340 34474 41368 35770
rect 41328 34468 41380 34474
rect 41328 34410 41380 34416
rect 40684 33992 40736 33998
rect 40684 33934 40736 33940
rect 41052 33992 41104 33998
rect 41052 33934 41104 33940
rect 40500 33924 40552 33930
rect 40500 33866 40552 33872
rect 40052 33782 40172 33810
rect 40052 32978 40080 33782
rect 40040 32972 40092 32978
rect 40040 32914 40092 32920
rect 40052 32434 40080 32914
rect 40316 32768 40368 32774
rect 40316 32710 40368 32716
rect 40040 32428 40092 32434
rect 40040 32370 40092 32376
rect 40040 32292 40092 32298
rect 40040 32234 40092 32240
rect 40052 31822 40080 32234
rect 40328 32026 40356 32710
rect 40408 32360 40460 32366
rect 40408 32302 40460 32308
rect 40316 32020 40368 32026
rect 40316 31962 40368 31968
rect 39396 31816 39448 31822
rect 39396 31758 39448 31764
rect 40040 31816 40092 31822
rect 40040 31758 40092 31764
rect 39212 31680 39264 31686
rect 39212 31622 39264 31628
rect 39224 31414 39252 31622
rect 40420 31482 40448 32302
rect 40408 31476 40460 31482
rect 40408 31418 40460 31424
rect 39212 31408 39264 31414
rect 39212 31350 39264 31356
rect 38936 31340 38988 31346
rect 38936 31282 38988 31288
rect 40040 30592 40092 30598
rect 40040 30534 40092 30540
rect 38844 30252 38896 30258
rect 38844 30194 38896 30200
rect 39764 30252 39816 30258
rect 39764 30194 39816 30200
rect 38856 29714 38884 30194
rect 38936 30048 38988 30054
rect 38936 29990 38988 29996
rect 38844 29708 38896 29714
rect 38844 29650 38896 29656
rect 38948 29646 38976 29990
rect 39776 29850 39804 30194
rect 40052 29850 40080 30534
rect 40512 30326 40540 33866
rect 40592 32292 40644 32298
rect 40592 32234 40644 32240
rect 40604 31822 40632 32234
rect 40592 31816 40644 31822
rect 40592 31758 40644 31764
rect 40592 31680 40644 31686
rect 40592 31622 40644 31628
rect 40604 31278 40632 31622
rect 40696 31346 40724 33934
rect 41432 33658 41460 37130
rect 42628 36922 42656 37130
rect 42616 36916 42668 36922
rect 42616 36858 42668 36864
rect 42800 36780 42852 36786
rect 42800 36722 42852 36728
rect 42812 35834 42840 36722
rect 43364 36106 43392 37198
rect 43352 36100 43404 36106
rect 43352 36042 43404 36048
rect 42800 35828 42852 35834
rect 42800 35770 42852 35776
rect 43260 35828 43312 35834
rect 43260 35770 43312 35776
rect 42892 35692 42944 35698
rect 42892 35634 42944 35640
rect 42904 35290 42932 35634
rect 42892 35284 42944 35290
rect 42892 35226 42944 35232
rect 43168 35080 43220 35086
rect 43168 35022 43220 35028
rect 42800 35012 42852 35018
rect 42800 34954 42852 34960
rect 41420 33652 41472 33658
rect 41420 33594 41472 33600
rect 41236 33584 41288 33590
rect 41236 33526 41288 33532
rect 40868 33516 40920 33522
rect 40868 33458 40920 33464
rect 40880 32842 40908 33458
rect 41052 33380 41104 33386
rect 41052 33322 41104 33328
rect 41064 32978 41092 33322
rect 41144 33312 41196 33318
rect 41144 33254 41196 33260
rect 41052 32972 41104 32978
rect 41052 32914 41104 32920
rect 40868 32836 40920 32842
rect 40868 32778 40920 32784
rect 40880 32450 40908 32778
rect 41064 32502 41092 32914
rect 40788 32422 40908 32450
rect 41052 32496 41104 32502
rect 41052 32438 41104 32444
rect 40788 31958 40816 32422
rect 40868 32360 40920 32366
rect 40868 32302 40920 32308
rect 40880 32026 40908 32302
rect 40960 32224 41012 32230
rect 40960 32166 41012 32172
rect 40868 32020 40920 32026
rect 40868 31962 40920 31968
rect 40776 31952 40828 31958
rect 40776 31894 40828 31900
rect 40788 31822 40816 31894
rect 40776 31816 40828 31822
rect 40776 31758 40828 31764
rect 40972 31754 41000 32166
rect 41064 31890 41092 32438
rect 41156 32434 41184 33254
rect 41248 32502 41276 33526
rect 42616 32972 42668 32978
rect 42616 32914 42668 32920
rect 41788 32836 41840 32842
rect 41788 32778 41840 32784
rect 41328 32768 41380 32774
rect 41328 32710 41380 32716
rect 41236 32496 41288 32502
rect 41236 32438 41288 32444
rect 41144 32428 41196 32434
rect 41144 32370 41196 32376
rect 41144 32224 41196 32230
rect 41144 32166 41196 32172
rect 41052 31884 41104 31890
rect 41052 31826 41104 31832
rect 40960 31748 41012 31754
rect 40960 31690 41012 31696
rect 40684 31340 40736 31346
rect 40684 31282 40736 31288
rect 41156 31278 41184 32166
rect 41248 31890 41276 32438
rect 41340 32314 41368 32710
rect 41800 32570 41828 32778
rect 41604 32564 41656 32570
rect 41604 32506 41656 32512
rect 41788 32564 41840 32570
rect 41788 32506 41840 32512
rect 41880 32564 41932 32570
rect 41880 32506 41932 32512
rect 41616 32473 41644 32506
rect 41602 32464 41658 32473
rect 41420 32428 41472 32434
rect 41602 32399 41658 32408
rect 41696 32428 41748 32434
rect 41420 32370 41472 32376
rect 41696 32370 41748 32376
rect 41432 32314 41460 32370
rect 41340 32286 41460 32314
rect 41236 31884 41288 31890
rect 41236 31826 41288 31832
rect 41340 31278 41368 32286
rect 41708 31770 41736 32370
rect 41892 32366 41920 32506
rect 42628 32434 42656 32914
rect 42616 32428 42668 32434
rect 42616 32370 42668 32376
rect 41880 32360 41932 32366
rect 42812 32314 42840 34954
rect 43180 33114 43208 35022
rect 43272 34610 43300 35770
rect 43364 35766 43392 36042
rect 43352 35760 43404 35766
rect 43352 35702 43404 35708
rect 43364 35222 43392 35702
rect 43352 35216 43404 35222
rect 43352 35158 43404 35164
rect 43260 34604 43312 34610
rect 43260 34546 43312 34552
rect 43168 33108 43220 33114
rect 43168 33050 43220 33056
rect 43180 32434 43208 33050
rect 43272 32570 43300 34546
rect 43364 32910 43392 35158
rect 43548 35086 43576 38830
rect 43720 38752 43772 38758
rect 43720 38694 43772 38700
rect 43732 38282 43760 38694
rect 43720 38276 43772 38282
rect 43720 38218 43772 38224
rect 44100 37262 44128 39986
rect 44744 39982 44772 40462
rect 45296 40186 45324 40462
rect 45284 40180 45336 40186
rect 45284 40122 45336 40128
rect 45008 40044 45060 40050
rect 45008 39986 45060 39992
rect 44180 39976 44232 39982
rect 44180 39918 44232 39924
rect 44732 39976 44784 39982
rect 44732 39918 44784 39924
rect 44192 38962 44220 39918
rect 44180 38956 44232 38962
rect 44180 38898 44232 38904
rect 44456 38956 44508 38962
rect 44456 38898 44508 38904
rect 44364 38888 44416 38894
rect 44364 38830 44416 38836
rect 44272 38752 44324 38758
rect 44272 38694 44324 38700
rect 44284 38350 44312 38694
rect 44376 38350 44404 38830
rect 44468 38486 44496 38898
rect 44548 38752 44600 38758
rect 44548 38694 44600 38700
rect 44456 38480 44508 38486
rect 44456 38422 44508 38428
rect 44272 38344 44324 38350
rect 44272 38286 44324 38292
rect 44364 38344 44416 38350
rect 44364 38286 44416 38292
rect 44284 38026 44312 38286
rect 44560 38214 44588 38694
rect 44744 38418 44772 39918
rect 45020 39642 45048 39986
rect 45008 39636 45060 39642
rect 45008 39578 45060 39584
rect 45296 38894 45324 40122
rect 45376 39840 45428 39846
rect 45376 39782 45428 39788
rect 45388 39438 45416 39782
rect 45376 39432 45428 39438
rect 45376 39374 45428 39380
rect 45560 38956 45612 38962
rect 45560 38898 45612 38904
rect 45284 38888 45336 38894
rect 45284 38830 45336 38836
rect 45468 38888 45520 38894
rect 45468 38830 45520 38836
rect 45100 38480 45152 38486
rect 45100 38422 45152 38428
rect 44732 38412 44784 38418
rect 44732 38354 44784 38360
rect 45112 38350 45140 38422
rect 45480 38418 45508 38830
rect 45572 38554 45600 38898
rect 45560 38548 45612 38554
rect 45560 38490 45612 38496
rect 45468 38412 45520 38418
rect 45468 38354 45520 38360
rect 45100 38344 45152 38350
rect 45100 38286 45152 38292
rect 45376 38344 45428 38350
rect 45376 38286 45428 38292
rect 44548 38208 44600 38214
rect 44548 38150 44600 38156
rect 44192 37998 44312 38026
rect 45112 38010 45140 38286
rect 45100 38004 45152 38010
rect 44192 37330 44220 37998
rect 45100 37946 45152 37952
rect 44272 37868 44324 37874
rect 44272 37810 44324 37816
rect 44180 37324 44232 37330
rect 44180 37266 44232 37272
rect 44284 37262 44312 37810
rect 44088 37256 44140 37262
rect 44088 37198 44140 37204
rect 44272 37256 44324 37262
rect 44272 37198 44324 37204
rect 45388 37194 45416 38286
rect 45376 37188 45428 37194
rect 45376 37130 45428 37136
rect 44180 36168 44232 36174
rect 44232 36128 44312 36156
rect 44180 36110 44232 36116
rect 43996 36100 44048 36106
rect 43996 36042 44048 36048
rect 43444 35080 43496 35086
rect 43444 35022 43496 35028
rect 43536 35080 43588 35086
rect 43536 35022 43588 35028
rect 43456 34746 43484 35022
rect 43444 34740 43496 34746
rect 43444 34682 43496 34688
rect 44008 34202 44036 36042
rect 44180 36032 44232 36038
rect 44180 35974 44232 35980
rect 44192 35086 44220 35974
rect 44284 35834 44312 36128
rect 44272 35828 44324 35834
rect 44272 35770 44324 35776
rect 44180 35080 44232 35086
rect 44180 35022 44232 35028
rect 44192 34746 44220 35022
rect 44180 34740 44232 34746
rect 44180 34682 44232 34688
rect 44284 34610 44312 35770
rect 45192 35692 45244 35698
rect 45192 35634 45244 35640
rect 44364 35624 44416 35630
rect 44364 35566 44416 35572
rect 44376 35494 44404 35566
rect 44364 35488 44416 35494
rect 44364 35430 44416 35436
rect 44272 34604 44324 34610
rect 44272 34546 44324 34552
rect 44376 34542 44404 35430
rect 45204 35154 45232 35634
rect 44548 35148 44600 35154
rect 44548 35090 44600 35096
rect 45192 35148 45244 35154
rect 45192 35090 45244 35096
rect 44560 34610 44588 35090
rect 44548 34604 44600 34610
rect 44548 34546 44600 34552
rect 44180 34536 44232 34542
rect 44180 34478 44232 34484
rect 44364 34536 44416 34542
rect 44364 34478 44416 34484
rect 43996 34196 44048 34202
rect 43996 34138 44048 34144
rect 44192 33998 44220 34478
rect 44180 33992 44232 33998
rect 44180 33934 44232 33940
rect 44180 33856 44232 33862
rect 44180 33798 44232 33804
rect 44192 33454 44220 33798
rect 44180 33448 44232 33454
rect 44180 33390 44232 33396
rect 44192 33046 44220 33390
rect 44560 33114 44588 34546
rect 45100 33516 45152 33522
rect 45100 33458 45152 33464
rect 44548 33108 44600 33114
rect 44548 33050 44600 33056
rect 44180 33040 44232 33046
rect 44180 32982 44232 32988
rect 43904 32972 43956 32978
rect 43904 32914 43956 32920
rect 43352 32904 43404 32910
rect 43352 32846 43404 32852
rect 43536 32904 43588 32910
rect 43536 32846 43588 32852
rect 43260 32564 43312 32570
rect 43260 32506 43312 32512
rect 43168 32428 43220 32434
rect 43168 32370 43220 32376
rect 41880 32302 41932 32308
rect 42720 32298 42840 32314
rect 42708 32292 42840 32298
rect 42760 32286 42840 32292
rect 42708 32234 42760 32240
rect 41616 31742 41736 31770
rect 41616 31346 41644 31742
rect 41604 31340 41656 31346
rect 41604 31282 41656 31288
rect 42812 31278 42840 32286
rect 43180 31958 43208 32370
rect 43168 31952 43220 31958
rect 43168 31894 43220 31900
rect 40592 31272 40644 31278
rect 40592 31214 40644 31220
rect 41144 31272 41196 31278
rect 41144 31214 41196 31220
rect 41328 31272 41380 31278
rect 41328 31214 41380 31220
rect 42800 31272 42852 31278
rect 42800 31214 42852 31220
rect 40604 30938 40632 31214
rect 40592 30932 40644 30938
rect 40592 30874 40644 30880
rect 40500 30320 40552 30326
rect 40500 30262 40552 30268
rect 40224 30252 40276 30258
rect 40224 30194 40276 30200
rect 39764 29844 39816 29850
rect 39764 29786 39816 29792
rect 40040 29844 40092 29850
rect 40040 29786 40092 29792
rect 40236 29646 40264 30194
rect 40512 29646 40540 30262
rect 40604 30258 40632 30874
rect 40776 30728 40828 30734
rect 40776 30670 40828 30676
rect 40788 30394 40816 30670
rect 41144 30660 41196 30666
rect 41144 30602 41196 30608
rect 41156 30394 41184 30602
rect 40776 30388 40828 30394
rect 40776 30330 40828 30336
rect 41144 30388 41196 30394
rect 41144 30330 41196 30336
rect 41340 30326 41368 31214
rect 42340 30796 42392 30802
rect 42340 30738 42392 30744
rect 41328 30320 41380 30326
rect 41328 30262 41380 30268
rect 40592 30252 40644 30258
rect 40592 30194 40644 30200
rect 40776 30252 40828 30258
rect 40776 30194 40828 30200
rect 40604 29646 40632 30194
rect 40788 29850 40816 30194
rect 40776 29844 40828 29850
rect 40776 29786 40828 29792
rect 38936 29640 38988 29646
rect 38936 29582 38988 29588
rect 40224 29640 40276 29646
rect 40224 29582 40276 29588
rect 40500 29640 40552 29646
rect 40500 29582 40552 29588
rect 40592 29640 40644 29646
rect 40592 29582 40644 29588
rect 38752 29232 38804 29238
rect 38752 29174 38804 29180
rect 38476 28960 38528 28966
rect 38476 28902 38528 28908
rect 38488 28150 38516 28902
rect 38476 28144 38528 28150
rect 38764 28098 38792 29174
rect 38948 29034 38976 29582
rect 40236 29306 40264 29582
rect 40788 29306 40816 29786
rect 41340 29714 41368 30262
rect 41972 30252 42024 30258
rect 41972 30194 42024 30200
rect 41328 29708 41380 29714
rect 41328 29650 41380 29656
rect 41984 29646 42012 30194
rect 41972 29640 42024 29646
rect 41972 29582 42024 29588
rect 41984 29306 42012 29582
rect 40224 29300 40276 29306
rect 40224 29242 40276 29248
rect 40776 29300 40828 29306
rect 40776 29242 40828 29248
rect 41972 29300 42024 29306
rect 41972 29242 42024 29248
rect 40684 29164 40736 29170
rect 40684 29106 40736 29112
rect 41512 29164 41564 29170
rect 41512 29106 41564 29112
rect 40224 29096 40276 29102
rect 40224 29038 40276 29044
rect 38936 29028 38988 29034
rect 38936 28970 38988 28976
rect 38948 28218 38976 28970
rect 39212 28688 39264 28694
rect 39212 28630 39264 28636
rect 38936 28212 38988 28218
rect 38936 28154 38988 28160
rect 38476 28086 38528 28092
rect 38488 28014 38516 28086
rect 38672 28070 38792 28098
rect 39120 28076 39172 28082
rect 38476 28008 38528 28014
rect 38476 27950 38528 27956
rect 38292 27056 38344 27062
rect 38292 26998 38344 27004
rect 38304 26790 38332 26998
rect 38292 26784 38344 26790
rect 38292 26726 38344 26732
rect 38488 26382 38516 27950
rect 38016 26376 38068 26382
rect 38016 26318 38068 26324
rect 38476 26376 38528 26382
rect 38476 26318 38528 26324
rect 37924 26240 37976 26246
rect 37924 26182 37976 26188
rect 37188 25900 37240 25906
rect 37188 25842 37240 25848
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 36912 25832 36964 25838
rect 36912 25774 36964 25780
rect 36924 25294 36952 25774
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 37096 25152 37148 25158
rect 37096 25094 37148 25100
rect 37740 25152 37792 25158
rect 37740 25094 37792 25100
rect 37108 24206 37136 25094
rect 37188 24744 37240 24750
rect 37188 24686 37240 24692
rect 37096 24200 37148 24206
rect 37096 24142 37148 24148
rect 36912 24064 36964 24070
rect 36912 24006 36964 24012
rect 36924 23118 36952 24006
rect 36912 23112 36964 23118
rect 36912 23054 36964 23060
rect 36820 22568 36872 22574
rect 36820 22510 36872 22516
rect 36726 19816 36782 19825
rect 36726 19751 36782 19760
rect 36832 19718 36860 22510
rect 37200 22012 37228 24686
rect 37752 24342 37780 25094
rect 37740 24336 37792 24342
rect 37740 24278 37792 24284
rect 37740 24200 37792 24206
rect 37740 24142 37792 24148
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 37292 23050 37320 24006
rect 37752 23866 37780 24142
rect 37740 23860 37792 23866
rect 37740 23802 37792 23808
rect 37648 23724 37700 23730
rect 37700 23684 37780 23712
rect 37648 23666 37700 23672
rect 37556 23520 37608 23526
rect 37608 23480 37688 23508
rect 37556 23462 37608 23468
rect 37660 23254 37688 23480
rect 37648 23248 37700 23254
rect 37648 23190 37700 23196
rect 37556 23112 37608 23118
rect 37556 23054 37608 23060
rect 37280 23044 37332 23050
rect 37280 22986 37332 22992
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37464 22976 37516 22982
rect 37464 22918 37516 22924
rect 37384 22710 37412 22918
rect 37476 22778 37504 22918
rect 37568 22778 37596 23054
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37556 22772 37608 22778
rect 37556 22714 37608 22720
rect 37372 22704 37424 22710
rect 37372 22646 37424 22652
rect 37280 22024 37332 22030
rect 37200 21984 37280 22012
rect 37280 21966 37332 21972
rect 37292 20466 37320 21966
rect 37660 21554 37688 23190
rect 37752 22642 37780 23684
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 37752 22506 37780 22578
rect 37740 22500 37792 22506
rect 37740 22442 37792 22448
rect 37752 21894 37780 22442
rect 37740 21888 37792 21894
rect 37740 21830 37792 21836
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 37752 21486 37780 21830
rect 37740 21480 37792 21486
rect 37740 21422 37792 21428
rect 37280 20460 37332 20466
rect 37280 20402 37332 20408
rect 37740 20256 37792 20262
rect 37844 20244 37872 25842
rect 37936 24342 37964 26182
rect 38028 24750 38056 26318
rect 38672 26246 38700 28070
rect 39120 28018 39172 28024
rect 39132 27674 39160 28018
rect 39120 27668 39172 27674
rect 39120 27610 39172 27616
rect 39224 27606 39252 28630
rect 40132 28620 40184 28626
rect 40132 28562 40184 28568
rect 40144 28218 40172 28562
rect 40236 28558 40264 29038
rect 40408 29028 40460 29034
rect 40408 28970 40460 28976
rect 40420 28558 40448 28970
rect 40696 28626 40724 29106
rect 40684 28620 40736 28626
rect 40684 28562 40736 28568
rect 41144 28620 41196 28626
rect 41144 28562 41196 28568
rect 40224 28552 40276 28558
rect 40224 28494 40276 28500
rect 40408 28552 40460 28558
rect 40408 28494 40460 28500
rect 40132 28212 40184 28218
rect 40132 28154 40184 28160
rect 39212 27600 39264 27606
rect 39212 27542 39264 27548
rect 40144 27402 40172 28154
rect 40236 27674 40264 28494
rect 40224 27668 40276 27674
rect 40224 27610 40276 27616
rect 40132 27396 40184 27402
rect 40132 27338 40184 27344
rect 39488 26580 39540 26586
rect 39488 26522 39540 26528
rect 39500 26382 39528 26522
rect 40236 26518 40264 27610
rect 40316 27600 40368 27606
rect 40316 27542 40368 27548
rect 40328 27470 40356 27542
rect 40316 27464 40368 27470
rect 40316 27406 40368 27412
rect 40420 27334 40448 28494
rect 41052 27396 41104 27402
rect 41052 27338 41104 27344
rect 40408 27328 40460 27334
rect 40408 27270 40460 27276
rect 40420 26586 40448 27270
rect 40408 26580 40460 26586
rect 40408 26522 40460 26528
rect 40224 26512 40276 26518
rect 40224 26454 40276 26460
rect 39488 26376 39540 26382
rect 39488 26318 39540 26324
rect 38752 26308 38804 26314
rect 38752 26250 38804 26256
rect 38660 26240 38712 26246
rect 38660 26182 38712 26188
rect 38200 25696 38252 25702
rect 38200 25638 38252 25644
rect 38016 24744 38068 24750
rect 38016 24686 38068 24692
rect 37924 24336 37976 24342
rect 37924 24278 37976 24284
rect 37936 23662 37964 24278
rect 37924 23656 37976 23662
rect 37924 23598 37976 23604
rect 38212 20534 38240 25638
rect 38764 25226 38792 26250
rect 40236 26246 40264 26454
rect 40132 26240 40184 26246
rect 40132 26182 40184 26188
rect 40224 26240 40276 26246
rect 40224 26182 40276 26188
rect 40144 25906 40172 26182
rect 40236 26042 40264 26182
rect 40224 26036 40276 26042
rect 40224 25978 40276 25984
rect 40132 25900 40184 25906
rect 40132 25842 40184 25848
rect 38844 25424 38896 25430
rect 38844 25366 38896 25372
rect 38752 25220 38804 25226
rect 38752 25162 38804 25168
rect 38764 24954 38792 25162
rect 38752 24948 38804 24954
rect 38752 24890 38804 24896
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 38764 24410 38792 24754
rect 38752 24404 38804 24410
rect 38752 24346 38804 24352
rect 38660 24268 38712 24274
rect 38660 24210 38712 24216
rect 38292 23520 38344 23526
rect 38672 23474 38700 24210
rect 38856 24206 38884 25366
rect 39028 25288 39080 25294
rect 39028 25230 39080 25236
rect 39040 24274 39068 25230
rect 39120 25152 39172 25158
rect 39120 25094 39172 25100
rect 39132 24954 39160 25094
rect 39120 24948 39172 24954
rect 39120 24890 39172 24896
rect 39028 24268 39080 24274
rect 39028 24210 39080 24216
rect 39132 24206 39160 24890
rect 40132 24268 40184 24274
rect 40132 24210 40184 24216
rect 38844 24200 38896 24206
rect 38844 24142 38896 24148
rect 39120 24200 39172 24206
rect 39120 24142 39172 24148
rect 39132 23526 39160 24142
rect 40144 23866 40172 24210
rect 40132 23860 40184 23866
rect 40132 23802 40184 23808
rect 40776 23860 40828 23866
rect 40776 23802 40828 23808
rect 39948 23792 40000 23798
rect 39948 23734 40000 23740
rect 39488 23588 39540 23594
rect 39488 23530 39540 23536
rect 38292 23462 38344 23468
rect 38304 23118 38332 23462
rect 38488 23446 38700 23474
rect 39120 23520 39172 23526
rect 39120 23462 39172 23468
rect 38488 23118 38516 23446
rect 38292 23112 38344 23118
rect 38292 23054 38344 23060
rect 38476 23112 38528 23118
rect 38476 23054 38528 23060
rect 38384 22976 38436 22982
rect 38384 22918 38436 22924
rect 38396 21962 38424 22918
rect 38384 21956 38436 21962
rect 38384 21898 38436 21904
rect 38488 21690 38516 23054
rect 39132 22658 39160 23462
rect 39304 23044 39356 23050
rect 39304 22986 39356 22992
rect 38856 22642 39160 22658
rect 39316 22642 39344 22986
rect 39500 22642 39528 23530
rect 39960 23050 39988 23734
rect 40040 23724 40092 23730
rect 40040 23666 40092 23672
rect 39948 23044 40000 23050
rect 39948 22986 40000 22992
rect 40052 22778 40080 23666
rect 40144 23118 40172 23802
rect 40224 23520 40276 23526
rect 40224 23462 40276 23468
rect 40132 23112 40184 23118
rect 40132 23054 40184 23060
rect 40236 23050 40264 23462
rect 40788 23118 40816 23802
rect 41064 23118 41092 27338
rect 41156 24750 41184 28562
rect 41524 28558 41552 29106
rect 42352 29102 42380 30738
rect 43272 30598 43300 32506
rect 43548 32366 43576 32846
rect 43812 32428 43864 32434
rect 43812 32370 43864 32376
rect 43536 32360 43588 32366
rect 43536 32302 43588 32308
rect 43352 32224 43404 32230
rect 43352 32166 43404 32172
rect 43364 30870 43392 32166
rect 43824 32026 43852 32370
rect 43812 32020 43864 32026
rect 43812 31962 43864 31968
rect 43916 31822 43944 32914
rect 44548 32904 44600 32910
rect 44548 32846 44600 32852
rect 44088 32360 44140 32366
rect 44088 32302 44140 32308
rect 44100 31958 44128 32302
rect 44088 31952 44140 31958
rect 44088 31894 44140 31900
rect 43904 31816 43956 31822
rect 43904 31758 43956 31764
rect 43536 31272 43588 31278
rect 43536 31214 43588 31220
rect 43352 30864 43404 30870
rect 43352 30806 43404 30812
rect 43548 30734 43576 31214
rect 44100 30938 44128 31894
rect 44560 31754 44588 32846
rect 44824 32768 44876 32774
rect 44824 32710 44876 32716
rect 44836 32570 44864 32710
rect 44824 32564 44876 32570
rect 44824 32506 44876 32512
rect 45112 31890 45140 33458
rect 45204 33454 45232 35090
rect 45376 33992 45428 33998
rect 45376 33934 45428 33940
rect 45192 33448 45244 33454
rect 45192 33390 45244 33396
rect 45204 32502 45232 33390
rect 45284 33312 45336 33318
rect 45284 33254 45336 33260
rect 45296 32978 45324 33254
rect 45284 32972 45336 32978
rect 45284 32914 45336 32920
rect 45296 32570 45324 32914
rect 45284 32564 45336 32570
rect 45284 32506 45336 32512
rect 45192 32496 45244 32502
rect 45192 32438 45244 32444
rect 45100 31884 45152 31890
rect 45100 31826 45152 31832
rect 44548 31748 44600 31754
rect 44548 31690 44600 31696
rect 44088 30932 44140 30938
rect 44088 30874 44140 30880
rect 43536 30728 43588 30734
rect 43536 30670 43588 30676
rect 42892 30592 42944 30598
rect 42892 30534 42944 30540
rect 43260 30592 43312 30598
rect 43260 30534 43312 30540
rect 42904 30326 42932 30534
rect 42892 30320 42944 30326
rect 42892 30262 42944 30268
rect 43076 30252 43128 30258
rect 43076 30194 43128 30200
rect 42892 30184 42944 30190
rect 42892 30126 42944 30132
rect 42340 29096 42392 29102
rect 42340 29038 42392 29044
rect 41512 28552 41564 28558
rect 41512 28494 41564 28500
rect 41604 28552 41656 28558
rect 41604 28494 41656 28500
rect 42432 28552 42484 28558
rect 42432 28494 42484 28500
rect 41524 28218 41552 28494
rect 41512 28212 41564 28218
rect 41512 28154 41564 28160
rect 41524 27538 41552 28154
rect 41616 27674 41644 28494
rect 42340 28416 42392 28422
rect 42340 28358 42392 28364
rect 42352 28150 42380 28358
rect 42340 28144 42392 28150
rect 42340 28086 42392 28092
rect 42444 27674 42472 28494
rect 42904 28014 42932 30126
rect 43088 29306 43116 30194
rect 44100 30122 44128 30874
rect 45008 30252 45060 30258
rect 45008 30194 45060 30200
rect 44088 30116 44140 30122
rect 44088 30058 44140 30064
rect 43628 30048 43680 30054
rect 43628 29990 43680 29996
rect 43640 29646 43668 29990
rect 45020 29646 45048 30194
rect 45112 30190 45140 31826
rect 45204 31822 45232 32438
rect 45192 31816 45244 31822
rect 45192 31758 45244 31764
rect 45388 30734 45416 33934
rect 45652 32904 45704 32910
rect 45652 32846 45704 32852
rect 45664 32026 45692 32846
rect 45652 32020 45704 32026
rect 45652 31962 45704 31968
rect 45756 30818 45784 45526
rect 45940 45082 45968 45834
rect 46860 45422 46888 46271
rect 47044 46102 47072 49200
rect 47214 49056 47270 49065
rect 47214 48991 47270 49000
rect 47228 47122 47256 48991
rect 47216 47116 47268 47122
rect 47216 47058 47268 47064
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 48134 47016 48190 47025
rect 47032 46096 47084 46102
rect 47032 46038 47084 46044
rect 47584 45824 47636 45830
rect 47584 45766 47636 45772
rect 46848 45416 46900 45422
rect 46848 45358 46900 45364
rect 46480 45280 46532 45286
rect 46480 45222 46532 45228
rect 45928 45076 45980 45082
rect 45928 45018 45980 45024
rect 46492 44946 46520 45222
rect 46480 44940 46532 44946
rect 46480 44882 46532 44888
rect 46664 44804 46716 44810
rect 46664 44746 46716 44752
rect 46676 44538 46704 44746
rect 46664 44532 46716 44538
rect 46664 44474 46716 44480
rect 47216 44192 47268 44198
rect 47216 44134 47268 44140
rect 47308 44192 47360 44198
rect 47308 44134 47360 44140
rect 47228 43858 47256 44134
rect 47216 43852 47268 43858
rect 47216 43794 47268 43800
rect 47124 43716 47176 43722
rect 47124 43658 47176 43664
rect 47136 43450 47164 43658
rect 47124 43444 47176 43450
rect 47124 43386 47176 43392
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 47044 43217 47072 43250
rect 47030 43208 47086 43217
rect 47030 43143 47086 43152
rect 47320 42294 47348 44134
rect 47492 43308 47544 43314
rect 47492 43250 47544 43256
rect 47308 42288 47360 42294
rect 47308 42230 47360 42236
rect 46480 42016 46532 42022
rect 46480 41958 46532 41964
rect 46492 41682 46520 41958
rect 46480 41676 46532 41682
rect 46480 41618 46532 41624
rect 46480 40928 46532 40934
rect 46480 40870 46532 40876
rect 46492 40594 46520 40870
rect 46480 40588 46532 40594
rect 46480 40530 46532 40536
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46492 39506 46520 39782
rect 46480 39500 46532 39506
rect 46480 39442 46532 39448
rect 46112 38344 46164 38350
rect 46112 38286 46164 38292
rect 46124 38010 46152 38286
rect 46848 38276 46900 38282
rect 46848 38218 46900 38224
rect 46860 38010 46888 38218
rect 46112 38004 46164 38010
rect 46112 37946 46164 37952
rect 46848 38004 46900 38010
rect 46848 37946 46900 37952
rect 46296 37868 46348 37874
rect 46296 37810 46348 37816
rect 46756 37868 46808 37874
rect 46756 37810 46808 37816
rect 47308 37868 47360 37874
rect 47308 37810 47360 37816
rect 46308 37466 46336 37810
rect 46296 37460 46348 37466
rect 46296 37402 46348 37408
rect 46204 37392 46256 37398
rect 46204 37334 46256 37340
rect 45836 37120 45888 37126
rect 45836 37062 45888 37068
rect 45848 30938 45876 37062
rect 45928 35148 45980 35154
rect 45928 35090 45980 35096
rect 45940 34542 45968 35090
rect 46020 35080 46072 35086
rect 46020 35022 46072 35028
rect 46032 34610 46060 35022
rect 46020 34604 46072 34610
rect 46020 34546 46072 34552
rect 45928 34536 45980 34542
rect 45928 34478 45980 34484
rect 45836 30932 45888 30938
rect 45836 30874 45888 30880
rect 45560 30796 45612 30802
rect 45756 30790 45968 30818
rect 45560 30738 45612 30744
rect 45376 30728 45428 30734
rect 45376 30670 45428 30676
rect 45192 30592 45244 30598
rect 45192 30534 45244 30540
rect 45204 30190 45232 30534
rect 45388 30258 45416 30670
rect 45376 30252 45428 30258
rect 45376 30194 45428 30200
rect 45100 30184 45152 30190
rect 45100 30126 45152 30132
rect 45192 30184 45244 30190
rect 45192 30126 45244 30132
rect 43628 29640 43680 29646
rect 43628 29582 43680 29588
rect 43720 29640 43772 29646
rect 43720 29582 43772 29588
rect 43996 29640 44048 29646
rect 43996 29582 44048 29588
rect 45008 29640 45060 29646
rect 45008 29582 45060 29588
rect 43260 29504 43312 29510
rect 43260 29446 43312 29452
rect 43272 29306 43300 29446
rect 43732 29306 43760 29582
rect 43076 29300 43128 29306
rect 43076 29242 43128 29248
rect 43260 29300 43312 29306
rect 43260 29242 43312 29248
rect 43720 29300 43772 29306
rect 43720 29242 43772 29248
rect 43904 29164 43956 29170
rect 43904 29106 43956 29112
rect 43812 28552 43864 28558
rect 43812 28494 43864 28500
rect 43168 28076 43220 28082
rect 43168 28018 43220 28024
rect 42892 28008 42944 28014
rect 42892 27950 42944 27956
rect 41604 27668 41656 27674
rect 41604 27610 41656 27616
rect 42432 27668 42484 27674
rect 42432 27610 42484 27616
rect 41512 27532 41564 27538
rect 41512 27474 41564 27480
rect 41616 27470 41644 27610
rect 41604 27464 41656 27470
rect 41604 27406 41656 27412
rect 42444 27334 42472 27610
rect 42904 27606 42932 27950
rect 43180 27674 43208 28018
rect 43824 27878 43852 28494
rect 43812 27872 43864 27878
rect 43812 27814 43864 27820
rect 43168 27668 43220 27674
rect 43168 27610 43220 27616
rect 42892 27600 42944 27606
rect 42892 27542 42944 27548
rect 43260 27600 43312 27606
rect 43260 27542 43312 27548
rect 42432 27328 42484 27334
rect 42432 27270 42484 27276
rect 41604 26852 41656 26858
rect 41604 26794 41656 26800
rect 41420 25220 41472 25226
rect 41420 25162 41472 25168
rect 41328 24812 41380 24818
rect 41328 24754 41380 24760
rect 41144 24744 41196 24750
rect 41144 24686 41196 24692
rect 41156 24342 41184 24686
rect 41340 24614 41368 24754
rect 41328 24608 41380 24614
rect 41328 24550 41380 24556
rect 41144 24336 41196 24342
rect 41144 24278 41196 24284
rect 41144 24064 41196 24070
rect 41144 24006 41196 24012
rect 40776 23112 40828 23118
rect 40776 23054 40828 23060
rect 41052 23112 41104 23118
rect 41052 23054 41104 23060
rect 40224 23044 40276 23050
rect 40224 22986 40276 22992
rect 40776 22976 40828 22982
rect 40776 22918 40828 22924
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40788 22642 40816 22918
rect 38844 22636 39172 22642
rect 38896 22630 39120 22636
rect 38844 22578 38896 22584
rect 39120 22578 39172 22584
rect 39304 22636 39356 22642
rect 39304 22578 39356 22584
rect 39488 22636 39540 22642
rect 39488 22578 39540 22584
rect 40776 22636 40828 22642
rect 40776 22578 40828 22584
rect 39028 22568 39080 22574
rect 39028 22510 39080 22516
rect 38476 21684 38528 21690
rect 38476 21626 38528 21632
rect 38476 20596 38528 20602
rect 38476 20538 38528 20544
rect 38200 20528 38252 20534
rect 38200 20470 38252 20476
rect 38016 20460 38068 20466
rect 38016 20402 38068 20408
rect 37792 20216 37872 20244
rect 37740 20198 37792 20204
rect 38028 20058 38056 20402
rect 38108 20256 38160 20262
rect 38108 20198 38160 20204
rect 38016 20052 38068 20058
rect 38016 19994 38068 20000
rect 36820 19712 36872 19718
rect 36820 19654 36872 19660
rect 36544 18760 36596 18766
rect 36544 18702 36596 18708
rect 36832 18290 36860 19654
rect 38120 19514 38148 20198
rect 38212 19990 38240 20470
rect 38200 19984 38252 19990
rect 38200 19926 38252 19932
rect 38212 19718 38240 19926
rect 38488 19854 38516 20538
rect 39040 20058 39068 22510
rect 41156 22030 41184 24006
rect 41340 23866 41368 24550
rect 41328 23860 41380 23866
rect 41328 23802 41380 23808
rect 41236 23044 41288 23050
rect 41236 22986 41288 22992
rect 40500 22024 40552 22030
rect 40500 21966 40552 21972
rect 41144 22024 41196 22030
rect 41144 21966 41196 21972
rect 40512 20330 40540 21966
rect 40500 20324 40552 20330
rect 40500 20266 40552 20272
rect 39120 20256 39172 20262
rect 39120 20198 39172 20204
rect 40512 20210 40540 20266
rect 39028 20052 39080 20058
rect 39028 19994 39080 20000
rect 38292 19848 38344 19854
rect 38476 19848 38528 19854
rect 38292 19790 38344 19796
rect 38474 19816 38476 19825
rect 38528 19816 38530 19825
rect 38200 19712 38252 19718
rect 38200 19654 38252 19660
rect 38304 19514 38332 19790
rect 38474 19751 38530 19760
rect 38108 19508 38160 19514
rect 38108 19450 38160 19456
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 38752 19440 38804 19446
rect 38752 19382 38804 19388
rect 38568 19304 38620 19310
rect 38568 19246 38620 19252
rect 38580 18426 38608 19246
rect 38660 19236 38712 19242
rect 38660 19178 38712 19184
rect 38672 18766 38700 19178
rect 38764 18766 38792 19382
rect 38936 19372 38988 19378
rect 38936 19314 38988 19320
rect 38948 18970 38976 19314
rect 38936 18964 38988 18970
rect 38936 18906 38988 18912
rect 39040 18834 39068 19994
rect 39132 19922 39160 20198
rect 40512 20182 40724 20210
rect 40132 19984 40184 19990
rect 40132 19926 40184 19932
rect 39120 19916 39172 19922
rect 39120 19858 39172 19864
rect 39132 19378 39160 19858
rect 40144 19854 40172 19926
rect 39488 19848 39540 19854
rect 39488 19790 39540 19796
rect 40132 19848 40184 19854
rect 40132 19790 40184 19796
rect 39500 19378 39528 19790
rect 40040 19712 40092 19718
rect 40040 19654 40092 19660
rect 39948 19440 40000 19446
rect 39948 19382 40000 19388
rect 39120 19372 39172 19378
rect 39120 19314 39172 19320
rect 39488 19372 39540 19378
rect 39488 19314 39540 19320
rect 39500 18902 39528 19314
rect 39960 19174 39988 19382
rect 40052 19378 40080 19654
rect 40040 19372 40092 19378
rect 40040 19314 40092 19320
rect 39672 19168 39724 19174
rect 39672 19110 39724 19116
rect 39948 19168 40000 19174
rect 39948 19110 40000 19116
rect 39488 18896 39540 18902
rect 39488 18838 39540 18844
rect 39684 18834 39712 19110
rect 39028 18828 39080 18834
rect 39028 18770 39080 18776
rect 39672 18828 39724 18834
rect 39672 18770 39724 18776
rect 38660 18760 38712 18766
rect 38660 18702 38712 18708
rect 38752 18760 38804 18766
rect 38752 18702 38804 18708
rect 38672 18426 38700 18702
rect 38568 18420 38620 18426
rect 38568 18362 38620 18368
rect 38660 18420 38712 18426
rect 38660 18362 38712 18368
rect 38764 18290 38792 18702
rect 36820 18284 36872 18290
rect 36820 18226 36872 18232
rect 38752 18284 38804 18290
rect 38752 18226 38804 18232
rect 40144 18222 40172 19790
rect 40592 19780 40644 19786
rect 40592 19722 40644 19728
rect 40224 19304 40276 19310
rect 40224 19246 40276 19252
rect 40236 18766 40264 19246
rect 40604 18902 40632 19722
rect 40696 19378 40724 20182
rect 41248 19938 41276 22986
rect 41432 21486 41460 25162
rect 41512 23724 41564 23730
rect 41512 23666 41564 23672
rect 41524 23594 41552 23666
rect 41512 23588 41564 23594
rect 41512 23530 41564 23536
rect 41616 23118 41644 26794
rect 43272 25906 43300 27542
rect 43352 27464 43404 27470
rect 43352 27406 43404 27412
rect 43364 26858 43392 27406
rect 43720 27396 43772 27402
rect 43824 27384 43852 27814
rect 43916 27674 43944 29106
rect 44008 28762 44036 29582
rect 45112 29578 45140 30126
rect 45204 29850 45232 30126
rect 45572 30054 45600 30738
rect 45836 30728 45888 30734
rect 45836 30670 45888 30676
rect 45848 30258 45876 30670
rect 45836 30252 45888 30258
rect 45836 30194 45888 30200
rect 45560 30048 45612 30054
rect 45560 29990 45612 29996
rect 45192 29844 45244 29850
rect 45192 29786 45244 29792
rect 45744 29640 45796 29646
rect 45744 29582 45796 29588
rect 45100 29572 45152 29578
rect 45100 29514 45152 29520
rect 44088 29504 44140 29510
rect 44088 29446 44140 29452
rect 44100 29238 44128 29446
rect 44088 29232 44140 29238
rect 44088 29174 44140 29180
rect 45652 29164 45704 29170
rect 45652 29106 45704 29112
rect 45560 29096 45612 29102
rect 45560 29038 45612 29044
rect 43996 28756 44048 28762
rect 43996 28698 44048 28704
rect 43904 27668 43956 27674
rect 43904 27610 43956 27616
rect 43772 27356 43852 27384
rect 43720 27338 43772 27344
rect 43628 27328 43680 27334
rect 43628 27270 43680 27276
rect 43640 26994 43668 27270
rect 43732 27062 43760 27338
rect 43916 27130 43944 27610
rect 45572 27606 45600 29038
rect 45664 28762 45692 29106
rect 45652 28756 45704 28762
rect 45652 28698 45704 28704
rect 45756 28642 45784 29582
rect 45848 28966 45876 30194
rect 45836 28960 45888 28966
rect 45836 28902 45888 28908
rect 45664 28614 45784 28642
rect 45848 28626 45876 28902
rect 45940 28642 45968 30790
rect 46032 30598 46060 34546
rect 46020 30592 46072 30598
rect 46020 30534 46072 30540
rect 46032 30054 46060 30534
rect 46216 30190 46244 37334
rect 46480 36576 46532 36582
rect 46480 36518 46532 36524
rect 46492 36242 46520 36518
rect 46480 36236 46532 36242
rect 46480 36178 46532 36184
rect 46664 35692 46716 35698
rect 46664 35634 46716 35640
rect 46676 34746 46704 35634
rect 46664 34740 46716 34746
rect 46664 34682 46716 34688
rect 46664 32428 46716 32434
rect 46664 32370 46716 32376
rect 46480 32292 46532 32298
rect 46480 32234 46532 32240
rect 46492 31346 46520 32234
rect 46676 32026 46704 32370
rect 46664 32020 46716 32026
rect 46664 31962 46716 31968
rect 46676 31890 46704 31962
rect 46664 31884 46716 31890
rect 46664 31826 46716 31832
rect 46768 31754 46796 37810
rect 47124 35760 47176 35766
rect 47124 35702 47176 35708
rect 47032 35488 47084 35494
rect 47032 35430 47084 35436
rect 47044 35086 47072 35430
rect 46940 35080 46992 35086
rect 46940 35022 46992 35028
rect 47032 35080 47084 35086
rect 47032 35022 47084 35028
rect 46848 34944 46900 34950
rect 46848 34886 46900 34892
rect 46860 34610 46888 34886
rect 46848 34604 46900 34610
rect 46848 34546 46900 34552
rect 46952 31890 46980 35022
rect 47136 34406 47164 35702
rect 47216 35692 47268 35698
rect 47216 35634 47268 35640
rect 47228 34474 47256 35634
rect 47216 34468 47268 34474
rect 47216 34410 47268 34416
rect 47124 34400 47176 34406
rect 47124 34342 47176 34348
rect 47136 32434 47164 34342
rect 47124 32428 47176 32434
rect 47044 32388 47124 32416
rect 46940 31884 46992 31890
rect 46940 31826 46992 31832
rect 46676 31726 46796 31754
rect 46940 31748 46992 31754
rect 46480 31340 46532 31346
rect 46480 31282 46532 31288
rect 46204 30184 46256 30190
rect 46204 30126 46256 30132
rect 46020 30048 46072 30054
rect 46020 29990 46072 29996
rect 45836 28620 45888 28626
rect 45560 27600 45612 27606
rect 45560 27542 45612 27548
rect 43904 27124 43956 27130
rect 43904 27066 43956 27072
rect 43720 27056 43772 27062
rect 43720 26998 43772 27004
rect 43628 26988 43680 26994
rect 43628 26930 43680 26936
rect 43352 26852 43404 26858
rect 43352 26794 43404 26800
rect 43640 26586 43668 26930
rect 43628 26580 43680 26586
rect 43628 26522 43680 26528
rect 43916 26382 43944 27066
rect 45572 26994 45600 27542
rect 45664 27538 45692 28614
rect 45940 28614 46060 28642
rect 45836 28562 45888 28568
rect 45744 28552 45796 28558
rect 45744 28494 45796 28500
rect 45756 28218 45784 28494
rect 45744 28212 45796 28218
rect 45744 28154 45796 28160
rect 45848 28150 45876 28562
rect 45928 28552 45980 28558
rect 45928 28494 45980 28500
rect 45836 28144 45888 28150
rect 45836 28086 45888 28092
rect 45940 28082 45968 28494
rect 45744 28076 45796 28082
rect 45744 28018 45796 28024
rect 45928 28076 45980 28082
rect 45928 28018 45980 28024
rect 45652 27532 45704 27538
rect 45652 27474 45704 27480
rect 45756 27418 45784 28018
rect 45940 27674 45968 28018
rect 45928 27668 45980 27674
rect 45928 27610 45980 27616
rect 45664 27390 45784 27418
rect 45560 26988 45612 26994
rect 45560 26930 45612 26936
rect 45664 26790 45692 27390
rect 45652 26784 45704 26790
rect 45652 26726 45704 26732
rect 43904 26376 43956 26382
rect 43904 26318 43956 26324
rect 44548 26376 44600 26382
rect 44548 26318 44600 26324
rect 43536 26240 43588 26246
rect 43536 26182 43588 26188
rect 43548 25906 43576 26182
rect 44560 26042 44588 26318
rect 45664 26314 45692 26726
rect 45652 26308 45704 26314
rect 45652 26250 45704 26256
rect 44548 26036 44600 26042
rect 44548 25978 44600 25984
rect 43260 25900 43312 25906
rect 43260 25842 43312 25848
rect 43536 25900 43588 25906
rect 43536 25842 43588 25848
rect 42248 25424 42300 25430
rect 42248 25366 42300 25372
rect 42156 25288 42208 25294
rect 42156 25230 42208 25236
rect 41972 25220 42024 25226
rect 41972 25162 42024 25168
rect 41984 24614 42012 25162
rect 42064 25152 42116 25158
rect 42064 25094 42116 25100
rect 41972 24608 42024 24614
rect 41972 24550 42024 24556
rect 41984 24410 42012 24550
rect 41972 24404 42024 24410
rect 41972 24346 42024 24352
rect 42076 24274 42104 25094
rect 42168 24954 42196 25230
rect 42156 24948 42208 24954
rect 42156 24890 42208 24896
rect 42064 24268 42116 24274
rect 42064 24210 42116 24216
rect 41696 23724 41748 23730
rect 41696 23666 41748 23672
rect 41708 23186 41736 23666
rect 42076 23662 42104 24210
rect 42260 24206 42288 25366
rect 42892 25152 42944 25158
rect 42892 25094 42944 25100
rect 42904 24818 42932 25094
rect 43272 24886 43300 25842
rect 43260 24880 43312 24886
rect 43260 24822 43312 24828
rect 42708 24812 42760 24818
rect 42892 24812 42944 24818
rect 42760 24772 42840 24800
rect 42708 24754 42760 24760
rect 42248 24200 42300 24206
rect 42248 24142 42300 24148
rect 42812 23730 42840 24772
rect 42892 24754 42944 24760
rect 43272 24274 43300 24822
rect 45560 24676 45612 24682
rect 45560 24618 45612 24624
rect 43904 24608 43956 24614
rect 43904 24550 43956 24556
rect 43260 24268 43312 24274
rect 43260 24210 43312 24216
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42064 23656 42116 23662
rect 42064 23598 42116 23604
rect 41972 23588 42024 23594
rect 41972 23530 42024 23536
rect 41696 23180 41748 23186
rect 41696 23122 41748 23128
rect 41604 23112 41656 23118
rect 41604 23054 41656 23060
rect 41708 22778 41736 23122
rect 41696 22772 41748 22778
rect 41696 22714 41748 22720
rect 41604 22704 41656 22710
rect 41604 22646 41656 22652
rect 41512 22432 41564 22438
rect 41512 22374 41564 22380
rect 41524 22234 41552 22374
rect 41616 22234 41644 22646
rect 41512 22228 41564 22234
rect 41512 22170 41564 22176
rect 41604 22228 41656 22234
rect 41604 22170 41656 22176
rect 41616 22030 41644 22170
rect 41604 22024 41656 22030
rect 41604 21966 41656 21972
rect 41420 21480 41472 21486
rect 41420 21422 41472 21428
rect 41616 20534 41644 21966
rect 41788 21888 41840 21894
rect 41788 21830 41840 21836
rect 41800 21554 41828 21830
rect 41696 21548 41748 21554
rect 41696 21490 41748 21496
rect 41788 21548 41840 21554
rect 41788 21490 41840 21496
rect 41604 20528 41656 20534
rect 41604 20470 41656 20476
rect 41328 20460 41380 20466
rect 41328 20402 41380 20408
rect 41340 20058 41368 20402
rect 41328 20052 41380 20058
rect 41328 19994 41380 20000
rect 41248 19910 41368 19938
rect 41340 19854 41368 19910
rect 41236 19848 41288 19854
rect 41236 19790 41288 19796
rect 41328 19848 41380 19854
rect 41328 19790 41380 19796
rect 41248 19514 41276 19790
rect 41708 19718 41736 21490
rect 41880 20256 41932 20262
rect 41880 20198 41932 20204
rect 41892 19854 41920 20198
rect 41984 20058 42012 23530
rect 43272 23186 43300 24210
rect 43916 23730 43944 24550
rect 44180 24404 44232 24410
rect 44180 24346 44232 24352
rect 44088 23792 44140 23798
rect 44088 23734 44140 23740
rect 43904 23724 43956 23730
rect 43904 23666 43956 23672
rect 43812 23520 43864 23526
rect 43812 23462 43864 23468
rect 42708 23180 42760 23186
rect 42708 23122 42760 23128
rect 43260 23180 43312 23186
rect 43260 23122 43312 23128
rect 42720 22234 42748 23122
rect 43824 23118 43852 23462
rect 43916 23118 43944 23666
rect 44100 23186 44128 23734
rect 44192 23186 44220 24346
rect 45572 23905 45600 24618
rect 45664 24614 45692 26250
rect 46032 25430 46060 28614
rect 46480 28076 46532 28082
rect 46480 28018 46532 28024
rect 46388 27872 46440 27878
rect 46388 27814 46440 27820
rect 46400 27062 46428 27814
rect 46492 27674 46520 28018
rect 46480 27668 46532 27674
rect 46480 27610 46532 27616
rect 46388 27056 46440 27062
rect 46388 26998 46440 27004
rect 46020 25424 46072 25430
rect 46020 25366 46072 25372
rect 45928 25288 45980 25294
rect 45928 25230 45980 25236
rect 45940 24800 45968 25230
rect 46112 25220 46164 25226
rect 46112 25162 46164 25168
rect 46020 24812 46072 24818
rect 45940 24772 46020 24800
rect 46020 24754 46072 24760
rect 45652 24608 45704 24614
rect 45652 24550 45704 24556
rect 45652 24200 45704 24206
rect 45652 24142 45704 24148
rect 45558 23896 45614 23905
rect 45558 23831 45614 23840
rect 45376 23656 45428 23662
rect 45376 23598 45428 23604
rect 45560 23656 45612 23662
rect 45560 23598 45612 23604
rect 44088 23180 44140 23186
rect 44088 23122 44140 23128
rect 44180 23180 44232 23186
rect 44180 23122 44232 23128
rect 43812 23112 43864 23118
rect 43812 23054 43864 23060
rect 43904 23112 43956 23118
rect 44100 23066 44128 23122
rect 43904 23054 43956 23060
rect 44008 23038 44128 23066
rect 43352 22636 43404 22642
rect 43352 22578 43404 22584
rect 43364 22234 43392 22578
rect 44008 22506 44036 23038
rect 44088 22976 44140 22982
rect 44088 22918 44140 22924
rect 44100 22778 44128 22918
rect 44088 22772 44140 22778
rect 44088 22714 44140 22720
rect 43996 22500 44048 22506
rect 43996 22442 44048 22448
rect 42708 22228 42760 22234
rect 42708 22170 42760 22176
rect 43352 22228 43404 22234
rect 43352 22170 43404 22176
rect 42064 21956 42116 21962
rect 42064 21898 42116 21904
rect 42076 21622 42104 21898
rect 42064 21616 42116 21622
rect 42064 21558 42116 21564
rect 42720 21010 42748 22170
rect 43996 22092 44048 22098
rect 43996 22034 44048 22040
rect 42708 21004 42760 21010
rect 42708 20946 42760 20952
rect 42984 20868 43036 20874
rect 42984 20810 43036 20816
rect 42996 20602 43024 20810
rect 42984 20596 43036 20602
rect 42984 20538 43036 20544
rect 43444 20460 43496 20466
rect 44008 20448 44036 22034
rect 44100 22030 44128 22714
rect 44192 22710 44220 23122
rect 44272 23044 44324 23050
rect 44272 22986 44324 22992
rect 44180 22704 44232 22710
rect 44180 22646 44232 22652
rect 44284 22574 44312 22986
rect 44456 22976 44508 22982
rect 44456 22918 44508 22924
rect 44468 22642 44496 22918
rect 45388 22710 45416 23598
rect 45572 23322 45600 23598
rect 45560 23316 45612 23322
rect 45560 23258 45612 23264
rect 45664 23118 45692 24142
rect 45652 23112 45704 23118
rect 45652 23054 45704 23060
rect 45376 22704 45428 22710
rect 45376 22646 45428 22652
rect 44456 22636 44508 22642
rect 44456 22578 44508 22584
rect 45100 22636 45152 22642
rect 45100 22578 45152 22584
rect 44272 22568 44324 22574
rect 44272 22510 44324 22516
rect 44088 22024 44140 22030
rect 44088 21966 44140 21972
rect 44180 21888 44232 21894
rect 44180 21830 44232 21836
rect 44192 21486 44220 21830
rect 44272 21548 44324 21554
rect 44272 21490 44324 21496
rect 44180 21480 44232 21486
rect 44180 21422 44232 21428
rect 44088 20460 44140 20466
rect 44008 20420 44088 20448
rect 43444 20402 43496 20408
rect 44088 20402 44140 20408
rect 43352 20324 43404 20330
rect 43352 20266 43404 20272
rect 41972 20052 42024 20058
rect 41972 19994 42024 20000
rect 41880 19848 41932 19854
rect 41880 19790 41932 19796
rect 41696 19712 41748 19718
rect 41696 19654 41748 19660
rect 41236 19508 41288 19514
rect 41236 19450 41288 19456
rect 41892 19378 41920 19790
rect 40684 19372 40736 19378
rect 40684 19314 40736 19320
rect 41880 19372 41932 19378
rect 41880 19314 41932 19320
rect 40592 18896 40644 18902
rect 40592 18838 40644 18844
rect 40224 18760 40276 18766
rect 40224 18702 40276 18708
rect 40236 18426 40264 18702
rect 40224 18420 40276 18426
rect 40224 18362 40276 18368
rect 41984 18290 42012 19994
rect 43364 19854 43392 20266
rect 43456 20058 43484 20402
rect 43996 20256 44048 20262
rect 43996 20198 44048 20204
rect 43444 20052 43496 20058
rect 43444 19994 43496 20000
rect 43168 19848 43220 19854
rect 43168 19790 43220 19796
rect 43352 19848 43404 19854
rect 43352 19790 43404 19796
rect 43180 19514 43208 19790
rect 43168 19508 43220 19514
rect 43168 19450 43220 19456
rect 43812 19508 43864 19514
rect 43812 19450 43864 19456
rect 43824 19378 43852 19450
rect 43812 19372 43864 19378
rect 43812 19314 43864 19320
rect 43824 18970 43852 19314
rect 43812 18964 43864 18970
rect 43812 18906 43864 18912
rect 44008 18766 44036 20198
rect 44100 19854 44128 20402
rect 44088 19848 44140 19854
rect 44088 19790 44140 19796
rect 44284 19310 44312 21490
rect 45112 21146 45140 22578
rect 45664 22438 45692 23054
rect 45652 22432 45704 22438
rect 45652 22374 45704 22380
rect 44640 21140 44692 21146
rect 44640 21082 44692 21088
rect 45100 21140 45152 21146
rect 45100 21082 45152 21088
rect 44652 20466 44680 21082
rect 44640 20460 44692 20466
rect 44640 20402 44692 20408
rect 44652 19922 44680 20402
rect 44640 19916 44692 19922
rect 44640 19858 44692 19864
rect 44364 19712 44416 19718
rect 44364 19654 44416 19660
rect 44376 19378 44404 19654
rect 44364 19372 44416 19378
rect 44364 19314 44416 19320
rect 45664 19334 45692 22374
rect 44272 19304 44324 19310
rect 44272 19246 44324 19252
rect 44376 18834 44404 19314
rect 45664 19306 45876 19334
rect 44364 18828 44416 18834
rect 44364 18770 44416 18776
rect 43996 18760 44048 18766
rect 43996 18702 44048 18708
rect 41972 18284 42024 18290
rect 41972 18226 42024 18232
rect 35624 18216 35676 18222
rect 35624 18158 35676 18164
rect 40132 18216 40184 18222
rect 40132 18158 40184 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 41420 10056 41472 10062
rect 41420 9998 41472 10004
rect 41432 9654 41460 9998
rect 41420 9648 41472 9654
rect 41420 9590 41472 9596
rect 45192 9648 45244 9654
rect 45192 9590 45244 9596
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 41432 8430 41460 9590
rect 44364 8492 44416 8498
rect 44364 8434 44416 8440
rect 41420 8424 41472 8430
rect 41420 8366 41472 8372
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24596 3738 24624 7346
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 44180 5024 44232 5030
rect 44180 4966 44232 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 40040 4616 40092 4622
rect 40040 4558 40092 4564
rect 38660 4072 38712 4078
rect 38660 4014 38712 4020
rect 39396 4072 39448 4078
rect 39396 4014 39448 4020
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24596 3534 24624 3674
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24780 3058 24808 3878
rect 25884 3602 25912 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 24964 3126 24992 3334
rect 24952 3120 25004 3126
rect 24952 3062 25004 3068
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 23860 800 23888 2382
rect 25792 800 25820 2926
rect 26436 800 26464 3538
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 27448 3058 27476 3470
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27540 2446 27568 3334
rect 31864 3058 31892 3470
rect 31852 3052 31904 3058
rect 31852 2994 31904 3000
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 27632 2650 27660 2926
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 27724 800 27752 2926
rect 32232 800 32260 2926
rect 32324 2446 32352 3470
rect 32496 3392 32548 3398
rect 32496 3334 32548 3340
rect 32508 3126 32536 3334
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 38396 3058 38424 3470
rect 38568 3392 38620 3398
rect 38568 3334 38620 3340
rect 38580 3126 38608 3334
rect 38568 3120 38620 3126
rect 38568 3062 38620 3068
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 38672 2650 38700 4014
rect 39304 4004 39356 4010
rect 39304 3946 39356 3952
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 39316 800 39344 3946
rect 39408 3602 39436 4014
rect 39396 3596 39448 3602
rect 39396 3538 39448 3544
rect 40052 2514 40080 4558
rect 40500 3936 40552 3942
rect 40500 3878 40552 3884
rect 42616 3936 42668 3942
rect 42616 3878 42668 3884
rect 42984 3936 43036 3942
rect 42984 3878 43036 3884
rect 40512 3602 40540 3878
rect 40500 3596 40552 3602
rect 40500 3538 40552 3544
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40224 2848 40276 2854
rect 40224 2790 40276 2796
rect 40236 2514 40264 2790
rect 40040 2508 40092 2514
rect 40040 2450 40092 2456
rect 40224 2508 40276 2514
rect 40224 2450 40276 2456
rect 40592 2508 40644 2514
rect 40592 2450 40644 2456
rect 40604 800 40632 2450
rect 41248 800 41276 3538
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 41420 3460 41472 3466
rect 41420 3402 41472 3408
rect 41432 3126 41460 3402
rect 41420 3120 41472 3126
rect 41420 3062 41472 3068
rect 42444 3058 42472 3470
rect 42628 3058 42656 3878
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 42812 3126 42840 3334
rect 42800 3120 42852 3126
rect 42800 3062 42852 3068
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 41880 2984 41932 2990
rect 41880 2926 41932 2932
rect 41892 800 41920 2926
rect 42996 2514 43024 3878
rect 44192 2582 44220 4966
rect 44272 4616 44324 4622
rect 44272 4558 44324 4564
rect 44284 3602 44312 4558
rect 44376 4146 44404 8434
rect 44548 5160 44600 5166
rect 44548 5102 44600 5108
rect 44560 4826 44588 5102
rect 44548 4820 44600 4826
rect 44548 4762 44600 4768
rect 45204 4622 45232 9590
rect 45848 6914 45876 19306
rect 46032 7886 46060 24754
rect 46124 24410 46152 25162
rect 46112 24404 46164 24410
rect 46112 24346 46164 24352
rect 46676 24206 46704 31726
rect 46940 31690 46992 31696
rect 46952 31210 46980 31690
rect 47044 31482 47072 32388
rect 47124 32370 47176 32376
rect 47124 32224 47176 32230
rect 47124 32166 47176 32172
rect 47136 31482 47164 32166
rect 47032 31476 47084 31482
rect 47032 31418 47084 31424
rect 47124 31476 47176 31482
rect 47124 31418 47176 31424
rect 46940 31204 46992 31210
rect 46940 31146 46992 31152
rect 47216 30048 47268 30054
rect 47216 29990 47268 29996
rect 47228 29714 47256 29990
rect 47216 29708 47268 29714
rect 47216 29650 47268 29656
rect 46848 28688 46900 28694
rect 46848 28630 46900 28636
rect 46860 27538 46888 28630
rect 46848 27532 46900 27538
rect 46848 27474 46900 27480
rect 46756 27464 46808 27470
rect 46756 27406 46808 27412
rect 46768 27130 46796 27406
rect 46756 27124 46808 27130
rect 46756 27066 46808 27072
rect 46940 26988 46992 26994
rect 46940 26930 46992 26936
rect 46848 25764 46900 25770
rect 46848 25706 46900 25712
rect 46860 24750 46888 25706
rect 46848 24744 46900 24750
rect 46848 24686 46900 24692
rect 46664 24200 46716 24206
rect 46664 24142 46716 24148
rect 46480 23112 46532 23118
rect 46480 23054 46532 23060
rect 46492 22710 46520 23054
rect 46480 22704 46532 22710
rect 46480 22646 46532 22652
rect 46480 22024 46532 22030
rect 46480 21966 46532 21972
rect 46492 21622 46520 21966
rect 46480 21616 46532 21622
rect 46480 21558 46532 21564
rect 46664 20256 46716 20262
rect 46664 20198 46716 20204
rect 46676 19922 46704 20198
rect 46664 19916 46716 19922
rect 46664 19858 46716 19864
rect 46480 17672 46532 17678
rect 46480 17614 46532 17620
rect 46492 17202 46520 17614
rect 46480 17196 46532 17202
rect 46480 17138 46532 17144
rect 46480 16992 46532 16998
rect 46480 16934 46532 16940
rect 46492 16658 46520 16934
rect 46480 16652 46532 16658
rect 46480 16594 46532 16600
rect 46664 14816 46716 14822
rect 46664 14758 46716 14764
rect 46676 14482 46704 14758
rect 46664 14476 46716 14482
rect 46664 14418 46716 14424
rect 46952 12850 46980 26930
rect 47216 25968 47268 25974
rect 47214 25936 47216 25945
rect 47268 25936 47270 25945
rect 47214 25871 47270 25880
rect 47124 25832 47176 25838
rect 47124 25774 47176 25780
rect 47136 24818 47164 25774
rect 47124 24812 47176 24818
rect 47124 24754 47176 24760
rect 47030 23488 47086 23497
rect 47030 23423 47086 23432
rect 47044 22642 47072 23423
rect 47124 23044 47176 23050
rect 47124 22986 47176 22992
rect 47136 22778 47164 22986
rect 47124 22772 47176 22778
rect 47124 22714 47176 22720
rect 47032 22636 47084 22642
rect 47032 22578 47084 22584
rect 47044 21554 47072 22578
rect 47124 21956 47176 21962
rect 47124 21898 47176 21904
rect 47136 21690 47164 21898
rect 47124 21684 47176 21690
rect 47124 21626 47176 21632
rect 47032 21548 47084 21554
rect 47032 21490 47084 21496
rect 47320 20466 47348 37810
rect 47400 37664 47452 37670
rect 47400 37606 47452 37612
rect 47412 34542 47440 37606
rect 47400 34536 47452 34542
rect 47400 34478 47452 34484
rect 47412 32366 47440 34478
rect 47400 32360 47452 32366
rect 47400 32302 47452 32308
rect 47400 32224 47452 32230
rect 47400 32166 47452 32172
rect 47412 24818 47440 32166
rect 47504 30258 47532 43250
rect 47492 30252 47544 30258
rect 47492 30194 47544 30200
rect 47492 28076 47544 28082
rect 47492 28018 47544 28024
rect 47400 24812 47452 24818
rect 47400 24754 47452 24760
rect 47032 20460 47084 20466
rect 47032 20402 47084 20408
rect 47308 20460 47360 20466
rect 47308 20402 47360 20408
rect 46940 12844 46992 12850
rect 46940 12786 46992 12792
rect 46846 12336 46902 12345
rect 46846 12271 46902 12280
rect 46664 11552 46716 11558
rect 46664 11494 46716 11500
rect 46676 11218 46704 11494
rect 46860 11218 46888 12271
rect 47044 11762 47072 20402
rect 47216 19372 47268 19378
rect 47216 19314 47268 19320
rect 47124 19168 47176 19174
rect 47124 19110 47176 19116
rect 47136 18834 47164 19110
rect 47124 18828 47176 18834
rect 47124 18770 47176 18776
rect 47124 13728 47176 13734
rect 47124 13670 47176 13676
rect 47136 13394 47164 13670
rect 47124 13388 47176 13394
rect 47124 13330 47176 13336
rect 47124 12640 47176 12646
rect 47124 12582 47176 12588
rect 47136 12306 47164 12582
rect 47124 12300 47176 12306
rect 47124 12242 47176 12248
rect 47032 11756 47084 11762
rect 47032 11698 47084 11704
rect 46664 11212 46716 11218
rect 46664 11154 46716 11160
rect 46848 11212 46900 11218
rect 46848 11154 46900 11160
rect 46020 7880 46072 7886
rect 46020 7822 46072 7828
rect 45756 6886 45876 6914
rect 45756 4622 45784 6886
rect 46480 6112 46532 6118
rect 46480 6054 46532 6060
rect 46664 6112 46716 6118
rect 46664 6054 46716 6060
rect 46020 5704 46072 5710
rect 46020 5646 46072 5652
rect 46032 5302 46060 5646
rect 46020 5296 46072 5302
rect 46020 5238 46072 5244
rect 45192 4616 45244 4622
rect 45192 4558 45244 4564
rect 45744 4616 45796 4622
rect 45744 4558 45796 4564
rect 45376 4480 45428 4486
rect 45376 4422 45428 4428
rect 44364 4140 44416 4146
rect 44364 4082 44416 4088
rect 44376 3738 44404 4082
rect 45100 3936 45152 3942
rect 45100 3878 45152 3884
rect 44364 3732 44416 3738
rect 44364 3674 44416 3680
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 44456 3528 44508 3534
rect 44456 3470 44508 3476
rect 44916 3528 44968 3534
rect 44916 3470 44968 3476
rect 44180 2576 44232 2582
rect 44180 2518 44232 2524
rect 44468 2514 44496 3470
rect 44928 3058 44956 3470
rect 45112 3126 45140 3878
rect 45100 3120 45152 3126
rect 45100 3062 45152 3068
rect 44916 3052 44968 3058
rect 44916 2994 44968 3000
rect 45100 2984 45152 2990
rect 45100 2926 45152 2932
rect 42984 2508 43036 2514
rect 42984 2450 43036 2456
rect 44456 2508 44508 2514
rect 44456 2450 44508 2456
rect 45112 800 45140 2926
rect 45388 2514 45416 4422
rect 45756 3194 45784 4558
rect 46492 4554 46520 6054
rect 46676 5778 46704 6054
rect 46664 5772 46716 5778
rect 46664 5714 46716 5720
rect 46480 4548 46532 4554
rect 46480 4490 46532 4496
rect 45836 4480 45888 4486
rect 45836 4422 45888 4428
rect 45848 3466 45876 4422
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 45836 3460 45888 3466
rect 45836 3402 45888 3408
rect 45744 3188 45796 3194
rect 45744 3130 45796 3136
rect 46756 2916 46808 2922
rect 46756 2858 46808 2864
rect 45376 2508 45428 2514
rect 45376 2450 45428 2456
rect 45744 2508 45796 2514
rect 45744 2450 45796 2456
rect 45756 800 45784 2450
rect 46768 1465 46796 2858
rect 46952 2650 46980 4014
rect 47044 3670 47072 11698
rect 47228 6322 47256 19314
rect 47504 18290 47532 28018
rect 47596 26994 47624 45766
rect 47688 44742 47716 46990
rect 47860 46980 47912 46986
rect 48134 46951 48190 46960
rect 47860 46922 47912 46928
rect 47872 45558 47900 46922
rect 48044 46504 48096 46510
rect 48044 46446 48096 46452
rect 48056 46170 48084 46446
rect 48044 46164 48096 46170
rect 48044 46106 48096 46112
rect 47860 45552 47912 45558
rect 47860 45494 47912 45500
rect 47676 44736 47728 44742
rect 47676 44678 47728 44684
rect 47688 37874 47716 44678
rect 47768 44396 47820 44402
rect 47768 44338 47820 44344
rect 47780 42226 47808 44338
rect 48148 43858 48176 46951
rect 48332 46646 48360 49200
rect 48320 46640 48372 46646
rect 48320 46582 48372 46588
rect 48226 44976 48282 44985
rect 48226 44911 48228 44920
rect 48280 44911 48282 44920
rect 48228 44882 48280 44888
rect 48320 44396 48372 44402
rect 48320 44338 48372 44344
rect 48136 43852 48188 43858
rect 48136 43794 48188 43800
rect 47860 43104 47912 43110
rect 47860 43046 47912 43052
rect 47872 42770 47900 43046
rect 48226 42936 48282 42945
rect 48226 42871 48282 42880
rect 48240 42770 48268 42871
rect 47860 42764 47912 42770
rect 47860 42706 47912 42712
rect 48228 42764 48280 42770
rect 48228 42706 48280 42712
rect 48332 42265 48360 44338
rect 48318 42256 48374 42265
rect 47768 42220 47820 42226
rect 48318 42191 48374 42200
rect 47768 42162 47820 42168
rect 47780 40050 47808 42162
rect 47860 42016 47912 42022
rect 47860 41958 47912 41964
rect 47872 41682 47900 41958
rect 47860 41676 47912 41682
rect 47860 41618 47912 41624
rect 48228 41676 48280 41682
rect 48228 41618 48280 41624
rect 48240 41585 48268 41618
rect 48226 41576 48282 41585
rect 48226 41511 48282 41520
rect 47860 40928 47912 40934
rect 47860 40870 47912 40876
rect 47872 40594 47900 40870
rect 47860 40588 47912 40594
rect 47860 40530 47912 40536
rect 48228 40588 48280 40594
rect 48228 40530 48280 40536
rect 48042 40216 48098 40225
rect 48042 40151 48098 40160
rect 47768 40044 47820 40050
rect 47768 39986 47820 39992
rect 47676 37868 47728 37874
rect 47676 37810 47728 37816
rect 47676 36848 47728 36854
rect 47676 36790 47728 36796
rect 47688 32230 47716 36790
rect 47676 32224 47728 32230
rect 47676 32166 47728 32172
rect 47676 30252 47728 30258
rect 47676 30194 47728 30200
rect 47584 26988 47636 26994
rect 47584 26930 47636 26936
rect 47688 19378 47716 30194
rect 47780 26330 47808 39986
rect 47860 39840 47912 39846
rect 47860 39782 47912 39788
rect 47872 39506 47900 39782
rect 47860 39500 47912 39506
rect 47860 39442 47912 39448
rect 47952 38752 48004 38758
rect 47952 38694 48004 38700
rect 47860 37664 47912 37670
rect 47860 37606 47912 37612
rect 47872 37194 47900 37606
rect 47860 37188 47912 37194
rect 47860 37130 47912 37136
rect 47964 37126 47992 38694
rect 48056 38418 48084 40151
rect 48240 39545 48268 40530
rect 48226 39536 48282 39545
rect 48136 39500 48188 39506
rect 48226 39471 48282 39480
rect 48136 39442 48188 39448
rect 48044 38412 48096 38418
rect 48044 38354 48096 38360
rect 48148 38185 48176 39442
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48226 37496 48282 37505
rect 48226 37431 48282 37440
rect 48240 37330 48268 37431
rect 48228 37324 48280 37330
rect 48228 37266 48280 37272
rect 47952 37120 48004 37126
rect 47952 37062 48004 37068
rect 47860 36576 47912 36582
rect 47860 36518 47912 36524
rect 47872 36242 47900 36518
rect 47860 36236 47912 36242
rect 47860 36178 47912 36184
rect 48228 36236 48280 36242
rect 48228 36178 48280 36184
rect 48240 36145 48268 36178
rect 48226 36136 48282 36145
rect 48226 36071 48282 36080
rect 48136 35556 48188 35562
rect 48136 35498 48188 35504
rect 48148 34202 48176 35498
rect 48136 34196 48188 34202
rect 48136 34138 48188 34144
rect 48320 33992 48372 33998
rect 48320 33934 48372 33940
rect 48332 33425 48360 33934
rect 48318 33416 48374 33425
rect 48318 33351 48374 33360
rect 47952 33312 48004 33318
rect 47952 33254 48004 33260
rect 47964 32978 47992 33254
rect 47952 32972 48004 32978
rect 47952 32914 48004 32920
rect 47860 32836 47912 32842
rect 47860 32778 47912 32784
rect 48320 32836 48372 32842
rect 48320 32778 48372 32784
rect 47872 32570 47900 32778
rect 48332 32745 48360 32778
rect 48318 32736 48374 32745
rect 48318 32671 48374 32680
rect 47860 32564 47912 32570
rect 47860 32506 47912 32512
rect 47858 32464 47914 32473
rect 47858 32399 47860 32408
rect 47912 32399 47914 32408
rect 48136 32428 48188 32434
rect 47860 32370 47912 32376
rect 48136 32370 48188 32376
rect 47860 30048 47912 30054
rect 47860 29990 47912 29996
rect 47872 29578 47900 29990
rect 47860 29572 47912 29578
rect 47860 29514 47912 29520
rect 47952 28960 48004 28966
rect 47952 28902 48004 28908
rect 47964 28626 47992 28902
rect 47952 28620 48004 28626
rect 47952 28562 48004 28568
rect 47860 28484 47912 28490
rect 47860 28426 47912 28432
rect 47872 28218 47900 28426
rect 47860 28212 47912 28218
rect 47860 28154 47912 28160
rect 47860 26784 47912 26790
rect 47860 26726 47912 26732
rect 47872 26450 47900 26726
rect 48042 26616 48098 26625
rect 48042 26551 48098 26560
rect 47860 26444 47912 26450
rect 47860 26386 47912 26392
rect 47780 26302 47900 26330
rect 47768 24812 47820 24818
rect 47768 24754 47820 24760
rect 47676 19372 47728 19378
rect 47676 19314 47728 19320
rect 47492 18284 47544 18290
rect 47492 18226 47544 18232
rect 47504 15026 47532 18226
rect 47780 16114 47808 24754
rect 47872 22094 47900 26302
rect 47952 26308 48004 26314
rect 47952 26250 48004 26256
rect 47964 25906 47992 26250
rect 47952 25900 48004 25906
rect 47952 25842 48004 25848
rect 48056 23798 48084 26551
rect 48044 23792 48096 23798
rect 48044 23734 48096 23740
rect 47872 22066 48084 22094
rect 47952 20256 48004 20262
rect 47952 20198 48004 20204
rect 47964 19990 47992 20198
rect 47952 19984 48004 19990
rect 47952 19926 48004 19932
rect 47952 19168 48004 19174
rect 47952 19110 48004 19116
rect 47964 18902 47992 19110
rect 47952 18896 48004 18902
rect 47952 18838 48004 18844
rect 47860 18080 47912 18086
rect 47860 18022 47912 18028
rect 47872 17746 47900 18022
rect 47860 17740 47912 17746
rect 47860 17682 47912 17688
rect 47860 16516 47912 16522
rect 47860 16458 47912 16464
rect 47872 16250 47900 16458
rect 47860 16244 47912 16250
rect 47860 16186 47912 16192
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47676 15496 47728 15502
rect 47676 15438 47728 15444
rect 47492 15020 47544 15026
rect 47492 14962 47544 14968
rect 47504 13938 47532 14962
rect 47688 14550 47716 15438
rect 47676 14544 47728 14550
rect 47676 14486 47728 14492
rect 47492 13932 47544 13938
rect 47492 13874 47544 13880
rect 47504 12434 47532 13874
rect 47504 12406 47624 12434
rect 47490 8256 47546 8265
rect 47490 8191 47546 8200
rect 47504 7954 47532 8191
rect 47492 7948 47544 7954
rect 47492 7890 47544 7896
rect 47596 6390 47624 12406
rect 47780 9654 47808 16050
rect 47952 13728 48004 13734
rect 47952 13670 48004 13676
rect 47964 13462 47992 13670
rect 47952 13456 48004 13462
rect 47952 13398 48004 13404
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 47964 12374 47992 12582
rect 47952 12368 48004 12374
rect 47952 12310 48004 12316
rect 47952 11552 48004 11558
rect 47952 11494 48004 11500
rect 47964 11286 47992 11494
rect 47952 11280 48004 11286
rect 47952 11222 48004 11228
rect 47768 9648 47820 9654
rect 47768 9590 47820 9596
rect 47952 7200 48004 7206
rect 47952 7142 48004 7148
rect 47964 6934 47992 7142
rect 47952 6928 48004 6934
rect 47952 6870 48004 6876
rect 47860 6724 47912 6730
rect 47860 6666 47912 6672
rect 47872 6458 47900 6666
rect 47860 6452 47912 6458
rect 47860 6394 47912 6400
rect 47584 6384 47636 6390
rect 47584 6326 47636 6332
rect 48056 6322 48084 22066
rect 47216 6316 47268 6322
rect 47216 6258 47268 6264
rect 47400 6316 47452 6322
rect 47400 6258 47452 6264
rect 48044 6316 48096 6322
rect 48044 6258 48096 6264
rect 47032 3664 47084 3670
rect 47032 3606 47084 3612
rect 47032 3460 47084 3466
rect 47032 3402 47084 3408
rect 46940 2644 46992 2650
rect 46940 2586 46992 2592
rect 46848 2304 46900 2310
rect 46848 2246 46900 2252
rect 46860 2145 46888 2246
rect 46846 2136 46902 2145
rect 46846 2071 46902 2080
rect 46754 1456 46810 1465
rect 46754 1391 46810 1400
rect 47044 800 47072 3402
rect 47412 3398 47440 6258
rect 47952 5636 48004 5642
rect 47952 5578 48004 5584
rect 47964 5234 47992 5578
rect 47952 5228 48004 5234
rect 47952 5170 48004 5176
rect 48148 4758 48176 32370
rect 48320 29572 48372 29578
rect 48320 29514 48372 29520
rect 48332 29345 48360 29514
rect 48318 29336 48374 29345
rect 48318 29271 48374 29280
rect 48226 28656 48282 28665
rect 48226 28591 48228 28600
rect 48280 28591 48282 28600
rect 48228 28562 48280 28568
rect 48226 27976 48282 27985
rect 48226 27911 48282 27920
rect 48240 26450 48268 27911
rect 48228 26444 48280 26450
rect 48228 26386 48280 26392
rect 48320 23044 48372 23050
rect 48320 22986 48372 22992
rect 48332 22545 48360 22986
rect 48318 22536 48374 22545
rect 48318 22471 48374 22480
rect 48320 21956 48372 21962
rect 48320 21898 48372 21904
rect 48332 21865 48360 21898
rect 48318 21856 48374 21865
rect 48318 21791 48374 21800
rect 48226 20496 48282 20505
rect 48226 20431 48282 20440
rect 48240 19922 48268 20431
rect 48228 19916 48280 19922
rect 48228 19858 48280 19864
rect 48226 19136 48282 19145
rect 48226 19071 48282 19080
rect 48240 18834 48268 19071
rect 48228 18828 48280 18834
rect 48228 18770 48280 18776
rect 48226 17776 48282 17785
rect 48226 17711 48228 17720
rect 48280 17711 48282 17720
rect 48228 17682 48280 17688
rect 48226 17096 48282 17105
rect 48226 17031 48282 17040
rect 48240 16658 48268 17031
rect 48228 16652 48280 16658
rect 48228 16594 48280 16600
rect 48226 15056 48282 15065
rect 48226 14991 48282 15000
rect 48240 14482 48268 14991
rect 48228 14476 48280 14482
rect 48228 14418 48280 14424
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 48240 13394 48268 13631
rect 48228 13388 48280 13394
rect 48228 13330 48280 13336
rect 48226 13016 48282 13025
rect 48226 12951 48282 12960
rect 48240 12306 48268 12951
rect 48228 12300 48280 12306
rect 48228 12242 48280 12248
rect 48226 6896 48282 6905
rect 48226 6831 48228 6840
rect 48280 6831 48282 6840
rect 48228 6802 48280 6808
rect 48228 5772 48280 5778
rect 48228 5714 48280 5720
rect 48240 5545 48268 5714
rect 48226 5536 48282 5545
rect 48226 5471 48282 5480
rect 48964 5160 49016 5166
rect 48964 5102 49016 5108
rect 48136 4752 48188 4758
rect 48136 4694 48188 4700
rect 47952 4684 48004 4690
rect 47952 4626 48004 4632
rect 47964 4146 47992 4626
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 47952 4140 48004 4146
rect 47952 4082 48004 4088
rect 47676 4072 47728 4078
rect 47676 4014 47728 4020
rect 47400 3392 47452 3398
rect 47400 3334 47452 3340
rect 47688 800 47716 4014
rect 47952 4004 48004 4010
rect 47952 3946 48004 3952
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47780 2446 47808 3878
rect 47964 3058 47992 3946
rect 47952 3052 48004 3058
rect 47952 2994 48004 3000
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 2566 200 2678 800
rect 3210 200 3322 800
rect 4498 200 4610 800
rect 5142 200 5254 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 15446 200 15558 800
rect 16090 200 16202 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 20598 200 20710 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25750 200 25862 800
rect 26394 200 26506 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 30258 200 30370 800
rect 30902 200 31014 800
rect 32190 200 32302 800
rect 32834 200 32946 800
rect 34122 200 34234 800
rect 34766 200 34878 800
rect 35410 200 35522 800
rect 36698 200 36810 800
rect 37342 200 37454 800
rect 38630 200 38742 800
rect 39274 200 39386 800
rect 40562 200 40674 800
rect 41206 200 41318 800
rect 41850 200 41962 800
rect 43138 200 43250 800
rect 43782 200 43894 800
rect 45070 200 45182 800
rect 45714 200 45826 800
rect 47002 200 47114 800
rect 47646 200 47758 800
rect 48332 105 48360 4490
rect 48976 800 49004 5102
rect 48934 200 49046 800
rect 49578 200 49690 800
rect 48318 96 48374 105
rect 48318 31 48374 40
<< via2 >>
rect 2778 48320 2834 48376
rect 3514 47640 3570 47696
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 2870 46280 2926 46336
rect 2778 45600 2834 45656
rect 2778 43560 2834 43616
rect 2778 40840 2834 40896
rect 2778 32680 2834 32736
rect 2778 25200 2834 25256
rect 2778 23840 2834 23896
rect 2778 21800 2834 21856
rect 2778 20440 2834 20496
rect 2778 18400 2834 18456
rect 2778 17076 2780 17096
rect 2780 17076 2832 17096
rect 2832 17076 2834 17096
rect 2778 17040 2834 17076
rect 2778 15000 2834 15056
rect 2778 14320 2834 14376
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 3514 41520 3570 41576
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 2962 10240 3018 10296
rect 2778 9560 2834 9616
rect 2962 7520 3018 7576
rect 2778 6840 2834 6896
rect 2962 5480 3018 5536
rect 2778 4800 2834 4856
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2962 3440 3018 3496
rect 2778 2760 2834 2816
rect 2870 1400 2926 1456
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 23846 27920 23902 27976
rect 24122 28076 24178 28112
rect 24122 28056 24124 28076
rect 24124 28056 24176 28076
rect 24176 28056 24178 28076
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 46846 46280 46902 46336
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 24766 28056 24822 28112
rect 25226 27940 25282 27976
rect 25226 27920 25228 27940
rect 25228 27920 25280 27940
rect 25280 27920 25282 27940
rect 27434 26832 27490 26888
rect 27894 26832 27950 26888
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 32770 20576 32826 20632
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34610 20576 34666 20632
rect 33506 20304 33562 20360
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 33966 19896 34022 19952
rect 35346 19896 35402 19952
rect 34610 19796 34612 19816
rect 34612 19796 34664 19816
rect 34664 19796 34666 19816
rect 34610 19760 34666 19796
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 36082 20304 36138 20360
rect 41602 32408 41658 32464
rect 36726 19760 36782 19816
rect 47214 49000 47270 49056
rect 47030 43152 47086 43208
rect 38474 19796 38476 19816
rect 38476 19796 38528 19816
rect 38528 19796 38530 19816
rect 38474 19760 38530 19796
rect 45558 23840 45614 23896
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 47214 25916 47216 25936
rect 47216 25916 47268 25936
rect 47268 25916 47270 25936
rect 47214 25880 47270 25916
rect 47030 23432 47086 23488
rect 46846 12280 46902 12336
rect 48134 46960 48190 47016
rect 48226 44940 48282 44976
rect 48226 44920 48228 44940
rect 48228 44920 48280 44940
rect 48280 44920 48282 44940
rect 48226 42880 48282 42936
rect 48318 42200 48374 42256
rect 48226 41520 48282 41576
rect 48042 40160 48098 40216
rect 48226 39480 48282 39536
rect 48134 38120 48190 38176
rect 48226 37440 48282 37496
rect 48226 36080 48282 36136
rect 48318 33360 48374 33416
rect 48318 32680 48374 32736
rect 47858 32428 47914 32464
rect 47858 32408 47860 32428
rect 47860 32408 47912 32428
rect 47912 32408 47914 32428
rect 48042 26560 48098 26616
rect 47490 8200 47546 8256
rect 46846 2080 46902 2136
rect 46754 1400 46810 1456
rect 48318 29280 48374 29336
rect 48226 28620 48282 28656
rect 48226 28600 48228 28620
rect 48228 28600 48280 28620
rect 48280 28600 48282 28620
rect 48226 27920 48282 27976
rect 48318 22480 48374 22536
rect 48318 21800 48374 21856
rect 48226 20440 48282 20496
rect 48226 19080 48282 19136
rect 48226 17740 48282 17776
rect 48226 17720 48228 17740
rect 48228 17720 48280 17740
rect 48280 17720 48282 17740
rect 48226 17040 48282 17096
rect 48226 15000 48282 15056
rect 48226 13640 48282 13696
rect 48226 12960 48282 13016
rect 48226 6860 48282 6896
rect 48226 6840 48228 6860
rect 48228 6840 48280 6860
rect 48280 6840 48282 6860
rect 48226 5480 48282 5536
rect 48318 40 48374 96
<< metal3 >>
rect 200 49588 800 49828
rect 47209 49058 47275 49061
rect 49200 49058 49800 49148
rect 47209 49056 49800 49058
rect 47209 49000 47214 49056
rect 47270 49000 49800 49056
rect 47209 48998 49800 49000
rect 47209 48995 47275 48998
rect 49200 48908 49800 48998
rect 200 48378 800 48468
rect 2773 48378 2839 48381
rect 200 48376 2839 48378
rect 200 48320 2778 48376
rect 2834 48320 2839 48376
rect 200 48318 2839 48320
rect 200 48228 800 48318
rect 2773 48315 2839 48318
rect 49200 48228 49800 48468
rect 200 47698 800 47788
rect 3509 47698 3575 47701
rect 200 47696 3575 47698
rect 200 47640 3514 47696
rect 3570 47640 3575 47696
rect 200 47638 3575 47640
rect 200 47548 800 47638
rect 3509 47635 3575 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 48129 47018 48195 47021
rect 49200 47018 49800 47108
rect 48129 47016 49800 47018
rect 48129 46960 48134 47016
rect 48190 46960 49800 47016
rect 48129 46958 49800 46960
rect 48129 46955 48195 46958
rect 49200 46868 49800 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 200 46338 800 46428
rect 2865 46338 2931 46341
rect 200 46336 2931 46338
rect 200 46280 2870 46336
rect 2926 46280 2931 46336
rect 200 46278 2931 46280
rect 200 46188 800 46278
rect 2865 46275 2931 46278
rect 46841 46338 46907 46341
rect 49200 46338 49800 46428
rect 46841 46336 49800 46338
rect 46841 46280 46846 46336
rect 46902 46280 49800 46336
rect 46841 46278 49800 46280
rect 46841 46275 46907 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 49200 46188 49800 46278
rect 200 45658 800 45748
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 2773 45658 2839 45661
rect 200 45656 2839 45658
rect 200 45600 2778 45656
rect 2834 45600 2839 45656
rect 200 45598 2839 45600
rect 200 45508 800 45598
rect 2773 45595 2839 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 48221 44978 48287 44981
rect 49200 44978 49800 45068
rect 48221 44976 49800 44978
rect 48221 44920 48226 44976
rect 48282 44920 49800 44976
rect 48221 44918 49800 44920
rect 48221 44915 48287 44918
rect 49200 44828 49800 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 200 44148 800 44388
rect 49200 44148 49800 44388
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 200 43618 800 43708
rect 2773 43618 2839 43621
rect 200 43616 2839 43618
rect 200 43560 2778 43616
rect 2834 43560 2839 43616
rect 200 43558 2839 43560
rect 200 43468 800 43558
rect 2773 43555 2839 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 47025 43210 47091 43213
rect 47158 43210 47164 43212
rect 47025 43208 47164 43210
rect 47025 43152 47030 43208
rect 47086 43152 47164 43208
rect 47025 43150 47164 43152
rect 47025 43147 47091 43150
rect 47158 43148 47164 43150
rect 47228 43148 47234 43212
rect 200 42788 800 43028
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 48221 42938 48287 42941
rect 49200 42938 49800 43028
rect 48221 42936 49800 42938
rect 48221 42880 48226 42936
rect 48282 42880 49800 42936
rect 48221 42878 49800 42880
rect 48221 42875 48287 42878
rect 49200 42788 49800 42878
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 48313 42258 48379 42261
rect 49200 42258 49800 42348
rect 48313 42256 49800 42258
rect 48313 42200 48318 42256
rect 48374 42200 49800 42256
rect 48313 42198 49800 42200
rect 48313 42195 48379 42198
rect 49200 42108 49800 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 200 41578 800 41668
rect 3509 41578 3575 41581
rect 200 41576 3575 41578
rect 200 41520 3514 41576
rect 3570 41520 3575 41576
rect 200 41518 3575 41520
rect 200 41428 800 41518
rect 3509 41515 3575 41518
rect 48221 41578 48287 41581
rect 49200 41578 49800 41668
rect 48221 41576 49800 41578
rect 48221 41520 48226 41576
rect 48282 41520 49800 41576
rect 48221 41518 49800 41520
rect 48221 41515 48287 41518
rect 49200 41428 49800 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 200 40898 800 40988
rect 2773 40898 2839 40901
rect 200 40896 2839 40898
rect 200 40840 2778 40896
rect 2834 40840 2839 40896
rect 200 40838 2839 40840
rect 200 40748 800 40838
rect 2773 40835 2839 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 48037 40218 48103 40221
rect 49200 40218 49800 40308
rect 48037 40216 49800 40218
rect 48037 40160 48042 40216
rect 48098 40160 49800 40216
rect 48037 40158 49800 40160
rect 48037 40155 48103 40158
rect 49200 40068 49800 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 200 39388 800 39628
rect 48221 39538 48287 39541
rect 49200 39538 49800 39628
rect 48221 39536 49800 39538
rect 48221 39480 48226 39536
rect 48282 39480 49800 39536
rect 48221 39478 49800 39480
rect 48221 39475 48287 39478
rect 49200 39388 49800 39478
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 200 38708 800 38948
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 48129 38178 48195 38181
rect 49200 38178 49800 38268
rect 48129 38176 49800 38178
rect 48129 38120 48134 38176
rect 48190 38120 49800 38176
rect 48129 38118 49800 38120
rect 48129 38115 48195 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 49200 38028 49800 38118
rect 200 37348 800 37588
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 48221 37498 48287 37501
rect 49200 37498 49800 37588
rect 48221 37496 49800 37498
rect 48221 37440 48226 37496
rect 48282 37440 49800 37496
rect 48221 37438 49800 37440
rect 48221 37435 48287 37438
rect 49200 37348 49800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36668 800 36908
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 35988 800 36228
rect 48221 36138 48287 36141
rect 49200 36138 49800 36228
rect 48221 36136 49800 36138
rect 48221 36080 48226 36136
rect 48282 36080 49800 36136
rect 48221 36078 49800 36080
rect 48221 36075 48287 36078
rect 49200 35988 49800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 49200 35308 49800 35548
rect 200 34628 800 34868
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 49200 34628 49800 34868
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 33948 800 34188
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 48313 33418 48379 33421
rect 49200 33418 49800 33508
rect 48313 33416 49800 33418
rect 48313 33360 48318 33416
rect 48374 33360 49800 33416
rect 48313 33358 49800 33360
rect 48313 33355 48379 33358
rect 49200 33268 49800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32828
rect 2773 32738 2839 32741
rect 200 32736 2839 32738
rect 200 32680 2778 32736
rect 2834 32680 2839 32736
rect 200 32678 2839 32680
rect 200 32588 800 32678
rect 2773 32675 2839 32678
rect 48313 32738 48379 32741
rect 49200 32738 49800 32828
rect 48313 32736 49800 32738
rect 48313 32680 48318 32736
rect 48374 32680 49800 32736
rect 48313 32678 49800 32680
rect 48313 32675 48379 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 49200 32588 49800 32678
rect 41597 32466 41663 32469
rect 47853 32466 47919 32469
rect 41597 32464 47919 32466
rect 41597 32408 41602 32464
rect 41658 32408 47858 32464
rect 47914 32408 47919 32464
rect 41597 32406 47919 32408
rect 41597 32403 41663 32406
rect 47853 32403 47919 32406
rect 200 31908 800 32148
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 49200 31228 49800 31468
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30548 800 30788
rect 49200 30548 49800 30788
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 200 29868 800 30108
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 200 29188 800 29428
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 48313 29338 48379 29341
rect 49200 29338 49800 29428
rect 48313 29336 49800 29338
rect 48313 29280 48318 29336
rect 48374 29280 49800 29336
rect 48313 29278 49800 29280
rect 48313 29275 48379 29278
rect 49200 29188 49800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 48221 28658 48287 28661
rect 49200 28658 49800 28748
rect 48221 28656 49800 28658
rect 48221 28600 48226 28656
rect 48282 28600 49800 28656
rect 48221 28598 49800 28600
rect 48221 28595 48287 28598
rect 49200 28508 49800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 24117 28114 24183 28117
rect 24761 28114 24827 28117
rect 24117 28112 24827 28114
rect 200 27828 800 28068
rect 24117 28056 24122 28112
rect 24178 28056 24766 28112
rect 24822 28056 24827 28112
rect 24117 28054 24827 28056
rect 24117 28051 24183 28054
rect 24761 28051 24827 28054
rect 23841 27978 23907 27981
rect 25221 27978 25287 27981
rect 23841 27976 25287 27978
rect 23841 27920 23846 27976
rect 23902 27920 25226 27976
rect 25282 27920 25287 27976
rect 23841 27918 25287 27920
rect 23841 27915 23907 27918
rect 25221 27915 25287 27918
rect 48221 27978 48287 27981
rect 49200 27978 49800 28068
rect 48221 27976 49800 27978
rect 48221 27920 48226 27976
rect 48282 27920 49800 27976
rect 48221 27918 49800 27920
rect 48221 27915 48287 27918
rect 49200 27828 49800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27148 800 27388
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 27429 26890 27495 26893
rect 27889 26890 27955 26893
rect 27429 26888 27955 26890
rect 27429 26832 27434 26888
rect 27490 26832 27894 26888
rect 27950 26832 27955 26888
rect 27429 26830 27955 26832
rect 27429 26827 27495 26830
rect 27889 26827 27955 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 48037 26618 48103 26621
rect 49200 26618 49800 26708
rect 48037 26616 49800 26618
rect 48037 26560 48042 26616
rect 48098 26560 49800 26616
rect 48037 26558 49800 26560
rect 48037 26555 48103 26558
rect 49200 26468 49800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25788 800 26028
rect 47209 25938 47275 25941
rect 49200 25938 49800 26028
rect 47209 25936 49800 25938
rect 47209 25880 47214 25936
rect 47270 25880 49800 25936
rect 47209 25878 49800 25880
rect 47209 25875 47275 25878
rect 49200 25788 49800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25348
rect 2773 25258 2839 25261
rect 200 25256 2839 25258
rect 200 25200 2778 25256
rect 2834 25200 2839 25256
rect 200 25198 2839 25200
rect 200 25108 800 25198
rect 2773 25195 2839 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 49200 24428 49800 24668
rect 200 23898 800 23988
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 2773 23898 2839 23901
rect 200 23896 2839 23898
rect 200 23840 2778 23896
rect 2834 23840 2839 23896
rect 200 23838 2839 23840
rect 200 23748 800 23838
rect 2773 23835 2839 23838
rect 45553 23898 45619 23901
rect 49200 23898 49800 23988
rect 45553 23896 49800 23898
rect 45553 23840 45558 23896
rect 45614 23840 49800 23896
rect 45553 23838 49800 23840
rect 45553 23835 45619 23838
rect 49200 23748 49800 23838
rect 47025 23490 47091 23493
rect 47158 23490 47164 23492
rect 47025 23488 47164 23490
rect 47025 23432 47030 23488
rect 47086 23432 47164 23488
rect 47025 23430 47164 23432
rect 47025 23427 47091 23430
rect 47158 23428 47164 23430
rect 47228 23428 47234 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23068 800 23308
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 48313 22538 48379 22541
rect 49200 22538 49800 22628
rect 48313 22536 49800 22538
rect 48313 22480 48318 22536
rect 48374 22480 49800 22536
rect 48313 22478 49800 22480
rect 48313 22475 48379 22478
rect 49200 22388 49800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 200 21858 800 21948
rect 2773 21858 2839 21861
rect 200 21856 2839 21858
rect 200 21800 2778 21856
rect 2834 21800 2839 21856
rect 200 21798 2839 21800
rect 200 21708 800 21798
rect 2773 21795 2839 21798
rect 48313 21858 48379 21861
rect 49200 21858 49800 21948
rect 48313 21856 49800 21858
rect 48313 21800 48318 21856
rect 48374 21800 49800 21856
rect 48313 21798 49800 21800
rect 48313 21795 48379 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 49200 21708 49800 21798
rect 200 21028 800 21268
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 32765 20634 32831 20637
rect 34605 20634 34671 20637
rect 32765 20632 34671 20634
rect 200 20498 800 20588
rect 32765 20576 32770 20632
rect 32826 20576 34610 20632
rect 34666 20576 34671 20632
rect 32765 20574 34671 20576
rect 32765 20571 32831 20574
rect 34605 20571 34671 20574
rect 2773 20498 2839 20501
rect 200 20496 2839 20498
rect 200 20440 2778 20496
rect 2834 20440 2839 20496
rect 200 20438 2839 20440
rect 200 20348 800 20438
rect 2773 20435 2839 20438
rect 48221 20498 48287 20501
rect 49200 20498 49800 20588
rect 48221 20496 49800 20498
rect 48221 20440 48226 20496
rect 48282 20440 49800 20496
rect 48221 20438 49800 20440
rect 48221 20435 48287 20438
rect 33501 20362 33567 20365
rect 36077 20362 36143 20365
rect 33501 20360 36143 20362
rect 33501 20304 33506 20360
rect 33562 20304 36082 20360
rect 36138 20304 36143 20360
rect 49200 20348 49800 20438
rect 33501 20302 36143 20304
rect 33501 20299 33567 20302
rect 36077 20299 36143 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 33961 19954 34027 19957
rect 35341 19954 35407 19957
rect 33961 19952 35407 19954
rect 33961 19896 33966 19952
rect 34022 19896 35346 19952
rect 35402 19896 35407 19952
rect 33961 19894 35407 19896
rect 33961 19891 34027 19894
rect 35341 19891 35407 19894
rect 34605 19818 34671 19821
rect 36721 19818 36787 19821
rect 38469 19818 38535 19821
rect 34605 19816 38535 19818
rect 34605 19760 34610 19816
rect 34666 19760 36726 19816
rect 36782 19760 38474 19816
rect 38530 19760 38535 19816
rect 34605 19758 38535 19760
rect 34605 19755 34671 19758
rect 36721 19755 36787 19758
rect 38469 19755 38535 19758
rect 49200 19668 49800 19908
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 18988 800 19228
rect 48221 19138 48287 19141
rect 49200 19138 49800 19228
rect 48221 19136 49800 19138
rect 48221 19080 48226 19136
rect 48282 19080 49800 19136
rect 48221 19078 49800 19080
rect 48221 19075 48287 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 49200 18988 49800 19078
rect 200 18458 800 18548
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 2773 18458 2839 18461
rect 200 18456 2839 18458
rect 200 18400 2778 18456
rect 2834 18400 2839 18456
rect 200 18398 2839 18400
rect 200 18308 800 18398
rect 2773 18395 2839 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 48221 17778 48287 17781
rect 49200 17778 49800 17868
rect 48221 17776 49800 17778
rect 48221 17720 48226 17776
rect 48282 17720 49800 17776
rect 48221 17718 49800 17720
rect 48221 17715 48287 17718
rect 49200 17628 49800 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 200 17098 800 17188
rect 2773 17098 2839 17101
rect 200 17096 2839 17098
rect 200 17040 2778 17096
rect 2834 17040 2839 17096
rect 200 17038 2839 17040
rect 200 16948 800 17038
rect 2773 17035 2839 17038
rect 48221 17098 48287 17101
rect 49200 17098 49800 17188
rect 48221 17096 49800 17098
rect 48221 17040 48226 17096
rect 48282 17040 49800 17096
rect 48221 17038 49800 17040
rect 48221 17035 48287 17038
rect 49200 16948 49800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 200 16268 800 16508
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 49200 15588 49800 15828
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 200 15058 800 15148
rect 2773 15058 2839 15061
rect 200 15056 2839 15058
rect 200 15000 2778 15056
rect 2834 15000 2839 15056
rect 200 14998 2839 15000
rect 200 14908 800 14998
rect 2773 14995 2839 14998
rect 48221 15058 48287 15061
rect 49200 15058 49800 15148
rect 48221 15056 49800 15058
rect 48221 15000 48226 15056
rect 48282 15000 49800 15056
rect 48221 14998 49800 15000
rect 48221 14995 48287 14998
rect 49200 14908 49800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14468
rect 2773 14378 2839 14381
rect 200 14376 2839 14378
rect 200 14320 2778 14376
rect 2834 14320 2839 14376
rect 200 14318 2839 14320
rect 200 14228 800 14318
rect 2773 14315 2839 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13548 800 13788
rect 48221 13698 48287 13701
rect 49200 13698 49800 13788
rect 48221 13696 49800 13698
rect 48221 13640 48226 13696
rect 48282 13640 49800 13696
rect 48221 13638 49800 13640
rect 48221 13635 48287 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 49200 13548 49800 13638
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 48221 13018 48287 13021
rect 49200 13018 49800 13108
rect 48221 13016 49800 13018
rect 48221 12960 48226 13016
rect 48282 12960 49800 13016
rect 48221 12958 49800 12960
rect 48221 12955 48287 12958
rect 49200 12868 49800 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12188 800 12428
rect 46841 12338 46907 12341
rect 49200 12338 49800 12428
rect 46841 12336 49800 12338
rect 46841 12280 46846 12336
rect 46902 12280 49800 12336
rect 46841 12278 49800 12280
rect 46841 12275 46907 12278
rect 49200 12188 49800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 200 11658 800 11748
rect 2773 11658 2839 11661
rect 200 11656 2839 11658
rect 200 11600 2778 11656
rect 2834 11600 2839 11656
rect 200 11598 2839 11600
rect 200 11508 800 11598
rect 2773 11595 2839 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 49200 10828 49800 11068
rect 200 10298 800 10388
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 2957 10298 3023 10301
rect 200 10296 3023 10298
rect 200 10240 2962 10296
rect 3018 10240 3023 10296
rect 200 10238 3023 10240
rect 200 10148 800 10238
rect 2957 10235 3023 10238
rect 49200 10148 49800 10388
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9708
rect 2773 9618 2839 9621
rect 200 9616 2839 9618
rect 200 9560 2778 9616
rect 2834 9560 2839 9616
rect 200 9558 2839 9560
rect 200 9468 800 9558
rect 2773 9555 2839 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 49200 8788 49800 9028
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 200 8108 800 8348
rect 47485 8258 47551 8261
rect 49200 8258 49800 8348
rect 47485 8256 49800 8258
rect 47485 8200 47490 8256
rect 47546 8200 49800 8256
rect 47485 8198 49800 8200
rect 47485 8195 47551 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 49200 8108 49800 8198
rect 200 7578 800 7668
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 2957 7578 3023 7581
rect 200 7576 3023 7578
rect 200 7520 2962 7576
rect 3018 7520 3023 7576
rect 200 7518 3023 7520
rect 200 7428 800 7518
rect 2957 7515 3023 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6988
rect 2773 6898 2839 6901
rect 200 6896 2839 6898
rect 200 6840 2778 6896
rect 2834 6840 2839 6896
rect 200 6838 2839 6840
rect 200 6748 800 6838
rect 2773 6835 2839 6838
rect 48221 6898 48287 6901
rect 49200 6898 49800 6988
rect 48221 6896 49800 6898
rect 48221 6840 48226 6896
rect 48282 6840 49800 6896
rect 48221 6838 49800 6840
rect 48221 6835 48287 6838
rect 49200 6748 49800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 49200 6068 49800 6308
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5628
rect 2957 5538 3023 5541
rect 200 5536 3023 5538
rect 200 5480 2962 5536
rect 3018 5480 3023 5536
rect 200 5478 3023 5480
rect 200 5388 800 5478
rect 2957 5475 3023 5478
rect 48221 5538 48287 5541
rect 49200 5538 49800 5628
rect 48221 5536 49800 5538
rect 48221 5480 48226 5536
rect 48282 5480 49800 5536
rect 48221 5478 49800 5480
rect 48221 5475 48287 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 49200 5388 49800 5478
rect 200 4858 800 4948
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 2773 4858 2839 4861
rect 200 4856 2839 4858
rect 200 4800 2778 4856
rect 2834 4800 2839 4856
rect 200 4798 2839 4800
rect 200 4708 800 4798
rect 2773 4795 2839 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 49200 4028 49800 4268
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3588
rect 2957 3498 3023 3501
rect 200 3496 3023 3498
rect 200 3440 2962 3496
rect 3018 3440 3023 3496
rect 200 3438 3023 3440
rect 200 3348 800 3438
rect 2957 3435 3023 3438
rect 49200 3348 49800 3588
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2908
rect 2773 2818 2839 2821
rect 200 2816 2839 2818
rect 200 2760 2778 2816
rect 2834 2760 2839 2816
rect 200 2758 2839 2760
rect 200 2668 800 2758
rect 2773 2755 2839 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 46841 2138 46907 2141
rect 49200 2138 49800 2228
rect 46841 2136 49800 2138
rect 46841 2080 46846 2136
rect 46902 2080 49800 2136
rect 46841 2078 49800 2080
rect 46841 2075 46907 2078
rect 49200 1988 49800 2078
rect 200 1458 800 1548
rect 2865 1458 2931 1461
rect 200 1456 2931 1458
rect 200 1400 2870 1456
rect 2926 1400 2931 1456
rect 200 1398 2931 1400
rect 200 1308 800 1398
rect 2865 1395 2931 1398
rect 46749 1458 46815 1461
rect 49200 1458 49800 1548
rect 46749 1456 49800 1458
rect 46749 1400 46754 1456
rect 46810 1400 49800 1456
rect 46749 1398 49800 1400
rect 46749 1395 46815 1398
rect 49200 1308 49800 1398
rect 200 628 800 868
rect 48313 98 48379 101
rect 49200 98 49800 188
rect 48313 96 49800 98
rect 48313 40 48318 96
rect 48374 40 49800 96
rect 48313 38 49800 40
rect 48313 35 48379 38
rect 49200 -52 49800 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 47164 43148 47228 43212
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 47164 23428 47228 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 47163 43212 47229 43213
rect 47163 43148 47164 43212
rect 47228 43148 47229 43212
rect 47163 43147 47229 43148
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 47166 23493 47226 43147
rect 47163 23492 47229 23493
rect 47163 23428 47164 23492
rect 47228 23428 47229 23492
rect 47163 23427 47229 23428
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform -1 0 24288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1667941163
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1667941163
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1667941163
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1667941163
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_290
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_302
timestamp 1667941163
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1667941163
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1667941163
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1667941163
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1667941163
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1667941163
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1667941163
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1667941163
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1667941163
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1667941163
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_510
timestamp 1667941163
transform 1 0 48024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1667941163
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1667941163
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_91
timestamp 1667941163
transform 1 0 9476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1667941163
transform 1 0 10212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1667941163
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1667941163
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_150
timestamp 1667941163
transform 1 0 14904 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1667941163
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_192
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_200
timestamp 1667941163
transform 1 0 19504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_248
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_256
timestamp 1667941163
transform 1 0 24656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1667941163
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_307
timestamp 1667941163
transform 1 0 29348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_319
timestamp 1667941163
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1667941163
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_360
timestamp 1667941163
transform 1 0 34224 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_372
timestamp 1667941163
transform 1 0 35328 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1667941163
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1667941163
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_440
timestamp 1667941163
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1667941163
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_472
timestamp 1667941163
transform 1 0 44528 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1667941163
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1667941163
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1667941163
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_510
timestamp 1667941163
transform 1 0 48024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1667941163
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1667941163
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1667941163
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1667941163
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1667941163
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1667941163
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_169
timestamp 1667941163
transform 1 0 16652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1667941163
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_180
timestamp 1667941163
transform 1 0 17664 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_188
timestamp 1667941163
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_216
timestamp 1667941163
transform 1 0 20976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_224
timestamp 1667941163
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_237
timestamp 1667941163
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1667941163
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1667941163
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_290
timestamp 1667941163
transform 1 0 27784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_297
timestamp 1667941163
transform 1 0 28428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1667941163
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_329
timestamp 1667941163
transform 1 0 31372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_342
timestamp 1667941163
transform 1 0 32568 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_354
timestamp 1667941163
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1667941163
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_404
timestamp 1667941163
transform 1 0 38272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_411
timestamp 1667941163
transform 1 0 38916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1667941163
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_421
timestamp 1667941163
transform 1 0 39836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_427
timestamp 1667941163
transform 1 0 40388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_449
timestamp 1667941163
transform 1 0 42412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_456
timestamp 1667941163
transform 1 0 43056 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_462
timestamp 1667941163
transform 1 0 43608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_466
timestamp 1667941163
transform 1 0 43976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1667941163
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_477
timestamp 1667941163
transform 1 0 44988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_483
timestamp 1667941163
transform 1 0 45540 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1667941163
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1667941163
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1667941163
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1667941163
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1667941163
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1667941163
transform 1 0 3404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1667941163
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 1667941163
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1667941163
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_74
timestamp 1667941163
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1667941163
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1667941163
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_128
timestamp 1667941163
transform 1 0 12880 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_132
timestamp 1667941163
transform 1 0 13248 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_144
timestamp 1667941163
transform 1 0 14352 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_156
timestamp 1667941163
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1667941163
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_269
timestamp 1667941163
transform 1 0 25852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_429
timestamp 1667941163
transform 1 0 40572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_436
timestamp 1667941163
transform 1 0 41216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_443
timestamp 1667941163
transform 1 0 41860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1667941163
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1667941163
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_461
timestamp 1667941163
transform 1 0 43516 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_466
timestamp 1667941163
transform 1 0 43976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_473
timestamp 1667941163
transform 1 0 44620 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1667941163
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1667941163
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_510
timestamp 1667941163
transform 1 0 48024 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_35
timestamp 1667941163
transform 1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1667941163
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_67
timestamp 1667941163
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1667941163
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1667941163
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1667941163
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_421
timestamp 1667941163
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_426
timestamp 1667941163
transform 1 0 40296 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_438
timestamp 1667941163
transform 1 0 41400 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_450
timestamp 1667941163
transform 1 0 42504 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_462
timestamp 1667941163
transform 1 0 43608 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_470
timestamp 1667941163
transform 1 0 44344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_474
timestamp 1667941163
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1667941163
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_482
timestamp 1667941163
transform 1 0 45448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_489
timestamp 1667941163
transform 1 0 46092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_514
timestamp 1667941163
transform 1 0 48392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1667941163
transform 1 0 4048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp 1667941163
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_47
timestamp 1667941163
transform 1 0 5428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1667941163
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1667941163
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1667941163
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1667941163
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1667941163
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1667941163
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1667941163
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_473
timestamp 1667941163
transform 1 0 44620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_477
timestamp 1667941163
transform 1 0 44988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1667941163
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_505
timestamp 1667941163
transform 1 0 47564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_510
timestamp 1667941163
transform 1 0 48024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1667941163
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1667941163
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1667941163
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_48
timestamp 1667941163
transform 1 0 5520 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_60
timestamp 1667941163
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_72
timestamp 1667941163
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1667941163
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1667941163
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1667941163
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1667941163
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1667941163
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1667941163
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1667941163
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1667941163
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_477
timestamp 1667941163
transform 1 0 44988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_485
timestamp 1667941163
transform 1 0 45724 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_489
timestamp 1667941163
transform 1 0 46092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_514
timestamp 1667941163
transform 1 0 48392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_32
timestamp 1667941163
transform 1 0 4048 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1667941163
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1667941163
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1667941163
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1667941163
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1667941163
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1667941163
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1667941163
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_485
timestamp 1667941163
transform 1 0 45724 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_491
timestamp 1667941163
transform 1 0 46276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_495
timestamp 1667941163
transform 1 0 46644 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_502
timestamp 1667941163
transform 1 0 47288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_505
timestamp 1667941163
transform 1 0 47564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_510
timestamp 1667941163
transform 1 0 48024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1667941163
transform 1 0 2392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1667941163
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_34
timestamp 1667941163
transform 1 0 4232 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_46
timestamp 1667941163
transform 1 0 5336 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_58
timestamp 1667941163
transform 1 0 6440 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_70
timestamp 1667941163
transform 1 0 7544 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1667941163
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1667941163
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1667941163
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1667941163
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1667941163
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1667941163
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1667941163
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1667941163
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1667941163
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_489
timestamp 1667941163
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_514
timestamp 1667941163
transform 1 0 48392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_31
timestamp 1667941163
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1667941163
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1667941163
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1667941163
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1667941163
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1667941163
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1667941163
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1667941163
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1667941163
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1667941163
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1667941163
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1667941163
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_505
timestamp 1667941163
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_510
timestamp 1667941163
transform 1 0 48024 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_46
timestamp 1667941163
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1667941163
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_70
timestamp 1667941163
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1667941163
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1667941163
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1667941163
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1667941163
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1667941163
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1667941163
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1667941163
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1667941163
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1667941163
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1667941163
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_501
timestamp 1667941163
transform 1 0 47196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_514
timestamp 1667941163
transform 1 0 48392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1667941163
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1667941163
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_429
timestamp 1667941163
transform 1 0 40572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_433
timestamp 1667941163
transform 1 0 40940 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1667941163
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1667941163
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1667941163
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1667941163
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1667941163
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1667941163
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1667941163
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1667941163
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1667941163
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1667941163
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1667941163
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1667941163
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1667941163
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1667941163
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1667941163
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1667941163
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1667941163
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1667941163
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1667941163
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1667941163
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1667941163
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1667941163
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1667941163
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1667941163
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1667941163
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1667941163
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1667941163
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1667941163
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1667941163
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1667941163
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1667941163
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1667941163
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1667941163
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1667941163
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1667941163
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1667941163
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1667941163
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1667941163
transform 1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1667941163
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1667941163
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1667941163
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1667941163
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1667941163
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1667941163
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1667941163
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1667941163
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1667941163
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1667941163
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1667941163
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1667941163
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1667941163
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1667941163
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1667941163
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1667941163
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1667941163
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1667941163
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1667941163
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1667941163
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1667941163
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1667941163
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1667941163
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1667941163
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1667941163
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1667941163
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1667941163
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1667941163
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1667941163
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1667941163
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1667941163
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1667941163
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1667941163
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1667941163
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1667941163
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_489
timestamp 1667941163
transform 1 0 46092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_514
timestamp 1667941163
transform 1 0 48392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_31
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_43
timestamp 1667941163
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1667941163
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1667941163
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1667941163
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1667941163
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1667941163
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1667941163
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1667941163
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1667941163
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_497
timestamp 1667941163
transform 1 0 46828 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_502
timestamp 1667941163
transform 1 0 47288 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_505
timestamp 1667941163
transform 1 0 47564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_510
timestamp 1667941163
transform 1 0 48024 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_14
timestamp 1667941163
transform 1 0 2392 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1667941163
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1667941163
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1667941163
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1667941163
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1667941163
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1667941163
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1667941163
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1667941163
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1667941163
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_489
timestamp 1667941163
transform 1 0 46092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_514
timestamp 1667941163
transform 1 0 48392 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1667941163
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1667941163
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1667941163
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1667941163
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1667941163
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1667941163
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1667941163
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1667941163
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_497
timestamp 1667941163
transform 1 0 46828 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1667941163
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_505
timestamp 1667941163
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_510
timestamp 1667941163
transform 1 0 48024 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1667941163
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1667941163
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1667941163
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1667941163
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1667941163
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1667941163
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1667941163
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1667941163
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1667941163
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_489
timestamp 1667941163
transform 1 0 46092 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_514
timestamp 1667941163
transform 1 0 48392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1667941163
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1667941163
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1667941163
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1667941163
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1667941163
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1667941163
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1667941163
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1667941163
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1667941163
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_497
timestamp 1667941163
transform 1 0 46828 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1667941163
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1667941163
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_510
timestamp 1667941163
transform 1 0 48024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1667941163
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1667941163
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1667941163
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1667941163
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1667941163
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1667941163
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1667941163
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1667941163
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1667941163
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_489
timestamp 1667941163
transform 1 0 46092 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_514
timestamp 1667941163
transform 1 0 48392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1667941163
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_31
timestamp 1667941163
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1667941163
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1667941163
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1667941163
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1667941163
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1667941163
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1667941163
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1667941163
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1667941163
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1667941163
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1667941163
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1667941163
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_505
timestamp 1667941163
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_510
timestamp 1667941163
transform 1 0 48024 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_10
timestamp 1667941163
transform 1 0 2024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_17
timestamp 1667941163
transform 1 0 2668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1667941163
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1667941163
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1667941163
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1667941163
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1667941163
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1667941163
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1667941163
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1667941163
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1667941163
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1667941163
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1667941163
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_501
timestamp 1667941163
transform 1 0 47196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_507
timestamp 1667941163
transform 1 0 47748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1667941163
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1667941163
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1667941163
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1667941163
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1667941163
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1667941163
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1667941163
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1667941163
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1667941163
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1667941163
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1667941163
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_505
timestamp 1667941163
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_510
timestamp 1667941163
transform 1 0 48024 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_14
timestamp 1667941163
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1667941163
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1667941163
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1667941163
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1667941163
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1667941163
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1667941163
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1667941163
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1667941163
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1667941163
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1667941163
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_489
timestamp 1667941163
transform 1 0 46092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_514
timestamp 1667941163
transform 1 0 48392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_31
timestamp 1667941163
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_43
timestamp 1667941163
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1667941163
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1667941163
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1667941163
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1667941163
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1667941163
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1667941163
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1667941163
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1667941163
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_497
timestamp 1667941163
transform 1 0 46828 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1667941163
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_505
timestamp 1667941163
transform 1 0 47564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_510
timestamp 1667941163
transform 1 0 48024 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1667941163
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1667941163
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1667941163
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1667941163
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1667941163
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1667941163
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1667941163
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1667941163
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1667941163
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1667941163
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_489
timestamp 1667941163
transform 1 0 46092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_514
timestamp 1667941163
transform 1 0 48392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1667941163
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_374
timestamp 1667941163
transform 1 0 35512 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1667941163
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_409
timestamp 1667941163
transform 1 0 38732 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_428
timestamp 1667941163
transform 1 0 40480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_440
timestamp 1667941163
transform 1 0 41584 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1667941163
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1667941163
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1667941163
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1667941163
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1667941163
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1667941163
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_505
timestamp 1667941163
transform 1 0 47564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_510
timestamp 1667941163
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_14
timestamp 1667941163
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1667941163
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1667941163
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_378
timestamp 1667941163
transform 1 0 35880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_390
timestamp 1667941163
transform 1 0 36984 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1667941163
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_412
timestamp 1667941163
transform 1 0 39008 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1667941163
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_430
timestamp 1667941163
transform 1 0 40664 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_442
timestamp 1667941163
transform 1 0 41768 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_454
timestamp 1667941163
transform 1 0 42872 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_462
timestamp 1667941163
transform 1 0 43608 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_467
timestamp 1667941163
transform 1 0 44068 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1667941163
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1667941163
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_489
timestamp 1667941163
transform 1 0 46092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_514
timestamp 1667941163
transform 1 0 48392 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1667941163
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_360
timestamp 1667941163
transform 1 0 34224 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_366
timestamp 1667941163
transform 1 0 34776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1667941163
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1667941163
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_399
timestamp 1667941163
transform 1 0 37812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_408
timestamp 1667941163
transform 1 0 38640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1667941163
transform 1 0 39744 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_431
timestamp 1667941163
transform 1 0 40756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_438
timestamp 1667941163
transform 1 0 41400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1667941163
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_449
timestamp 1667941163
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_464
timestamp 1667941163
transform 1 0 43792 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_474
timestamp 1667941163
transform 1 0 44712 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_486
timestamp 1667941163
transform 1 0 45816 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_498
timestamp 1667941163
transform 1 0 46920 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1667941163
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_505
timestamp 1667941163
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_510
timestamp 1667941163
transform 1 0 48024 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1667941163
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1667941163
transform 1 0 2668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1667941163
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_353
timestamp 1667941163
transform 1 0 33580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1667941163
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_373
timestamp 1667941163
transform 1 0 35420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_383
timestamp 1667941163
transform 1 0 36340 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_390
timestamp 1667941163
transform 1 0 36984 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_398
timestamp 1667941163
transform 1 0 37720 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_407
timestamp 1667941163
transform 1 0 38548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_414
timestamp 1667941163
transform 1 0 39192 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1667941163
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_429
timestamp 1667941163
transform 1 0 40572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_439
timestamp 1667941163
transform 1 0 41492 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_446
timestamp 1667941163
transform 1 0 42136 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_454
timestamp 1667941163
transform 1 0 42872 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_460
timestamp 1667941163
transform 1 0 43424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1667941163
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1667941163
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1667941163
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_489
timestamp 1667941163
transform 1 0 46092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_514
timestamp 1667941163
transform 1 0 48392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_9
timestamp 1667941163
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1667941163
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1667941163
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_243
timestamp 1667941163
transform 1 0 23460 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_255
timestamp 1667941163
transform 1 0 24564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1667941163
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_289
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_296
timestamp 1667941163
transform 1 0 28336 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_308
timestamp 1667941163
transform 1 0 29440 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1667941163
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_355
timestamp 1667941163
transform 1 0 33764 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_363
timestamp 1667941163
transform 1 0 34500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_380
timestamp 1667941163
transform 1 0 36064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_387
timestamp 1667941163
transform 1 0 36708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_397
timestamp 1667941163
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_414
timestamp 1667941163
transform 1 0 39192 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_426
timestamp 1667941163
transform 1 0 40296 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1667941163
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_449
timestamp 1667941163
transform 1 0 42412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_463
timestamp 1667941163
transform 1 0 43700 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_470
timestamp 1667941163
transform 1 0 44344 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_482
timestamp 1667941163
transform 1 0 45448 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_494
timestamp 1667941163
transform 1 0 46552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_498
timestamp 1667941163
transform 1 0 46920 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_502
timestamp 1667941163
transform 1 0 47288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_505
timestamp 1667941163
transform 1 0 47564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_510
timestamp 1667941163
transform 1 0 48024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_14
timestamp 1667941163
transform 1 0 2392 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1667941163
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_258
timestamp 1667941163
transform 1 0 24840 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_266
timestamp 1667941163
transform 1 0 25576 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_276
timestamp 1667941163
transform 1 0 26496 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_296
timestamp 1667941163
transform 1 0 28336 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_327
timestamp 1667941163
transform 1 0 31188 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_347
timestamp 1667941163
transform 1 0 33028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1667941163
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_383
timestamp 1667941163
transform 1 0 36340 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_395
timestamp 1667941163
transform 1 0 37444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_407
timestamp 1667941163
transform 1 0 38548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1667941163
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1667941163
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1667941163
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1667941163
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_457
timestamp 1667941163
transform 1 0 43148 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1667941163
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1667941163
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1667941163
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1667941163
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1667941163
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1667941163
transform 1 0 2392 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1667941163
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1667941163
transform 1 0 25852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1667941163
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_290
timestamp 1667941163
transform 1 0 27784 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_302
timestamp 1667941163
transform 1 0 28888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_310
timestamp 1667941163
transform 1 0 29624 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_316
timestamp 1667941163
transform 1 0 30176 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_328
timestamp 1667941163
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_400
timestamp 1667941163
transform 1 0 37904 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_412
timestamp 1667941163
transform 1 0 39008 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_424
timestamp 1667941163
transform 1 0 40112 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_436
timestamp 1667941163
transform 1 0 41216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1667941163
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1667941163
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_461
timestamp 1667941163
transform 1 0 43516 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_472
timestamp 1667941163
transform 1 0 44528 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_484
timestamp 1667941163
transform 1 0 45632 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_496
timestamp 1667941163
transform 1 0 46736 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1667941163
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1667941163
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_510
timestamp 1667941163
transform 1 0 48024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_327
timestamp 1667941163
transform 1 0 31188 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_339
timestamp 1667941163
transform 1 0 32292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_351
timestamp 1667941163
transform 1 0 33396 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_371
timestamp 1667941163
transform 1 0 35236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_383
timestamp 1667941163
transform 1 0 36340 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_391
timestamp 1667941163
transform 1 0 37076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_409
timestamp 1667941163
transform 1 0 38732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_417
timestamp 1667941163
transform 1 0 39468 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1667941163
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_436
timestamp 1667941163
transform 1 0 41216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_456
timestamp 1667941163
transform 1 0 43056 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_462
timestamp 1667941163
transform 1 0 43608 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_470
timestamp 1667941163
transform 1 0 44344 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1667941163
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_489
timestamp 1667941163
transform 1 0 46092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_514
timestamp 1667941163
transform 1 0 48392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_243
timestamp 1667941163
transform 1 0 23460 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_255
timestamp 1667941163
transform 1 0 24564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_267
timestamp 1667941163
transform 1 0 25668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1667941163
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_299
timestamp 1667941163
transform 1 0 28612 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_307
timestamp 1667941163
transform 1 0 29348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_314
timestamp 1667941163
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_322
timestamp 1667941163
transform 1 0 30728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_326
timestamp 1667941163
transform 1 0 31096 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1667941163
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_369
timestamp 1667941163
transform 1 0 35052 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1667941163
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_403
timestamp 1667941163
transform 1 0 38180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_420
timestamp 1667941163
transform 1 0 39744 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_440
timestamp 1667941163
transform 1 0 41584 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_449
timestamp 1667941163
transform 1 0 42412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_457
timestamp 1667941163
transform 1 0 43148 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_462
timestamp 1667941163
transform 1 0 43608 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_474
timestamp 1667941163
transform 1 0 44712 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_481
timestamp 1667941163
transform 1 0 45356 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_493
timestamp 1667941163
transform 1 0 46460 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1667941163
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_505
timestamp 1667941163
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_510
timestamp 1667941163
transform 1 0 48024 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_11
timestamp 1667941163
transform 1 0 2116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_17
timestamp 1667941163
transform 1 0 2668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1667941163
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_237
timestamp 1667941163
transform 1 0 22908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_272
timestamp 1667941163
transform 1 0 26128 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_280
timestamp 1667941163
transform 1 0 26864 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1667941163
transform 1 0 27600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 1667941163
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_317
timestamp 1667941163
transform 1 0 30268 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_324
timestamp 1667941163
transform 1 0 30912 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_344
timestamp 1667941163
transform 1 0 32752 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1667941163
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_372
timestamp 1667941163
transform 1 0 35328 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_390
timestamp 1667941163
transform 1 0 36984 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_400
timestamp 1667941163
transform 1 0 37904 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_407
timestamp 1667941163
transform 1 0 38548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1667941163
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1667941163
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_427
timestamp 1667941163
transform 1 0 40388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_435
timestamp 1667941163
transform 1 0 41124 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_439
timestamp 1667941163
transform 1 0 41492 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_460
timestamp 1667941163
transform 1 0 43424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_473
timestamp 1667941163
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_477
timestamp 1667941163
transform 1 0 44988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_483
timestamp 1667941163
transform 1 0 45540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_487
timestamp 1667941163
transform 1 0 45908 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_514
timestamp 1667941163
transform 1 0 48392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_31
timestamp 1667941163
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_43
timestamp 1667941163
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_235
timestamp 1667941163
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_246
timestamp 1667941163
transform 1 0 23736 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_258
timestamp 1667941163
transform 1 0 24840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_268
timestamp 1667941163
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_310
timestamp 1667941163
transform 1 0 29624 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_316
timestamp 1667941163
transform 1 0 30176 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_320
timestamp 1667941163
transform 1 0 30544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_353
timestamp 1667941163
transform 1 0 33580 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_357
timestamp 1667941163
transform 1 0 33948 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_369
timestamp 1667941163
transform 1 0 35052 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_377
timestamp 1667941163
transform 1 0 35788 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1667941163
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_399
timestamp 1667941163
transform 1 0 37812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_407
timestamp 1667941163
transform 1 0 38548 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_413
timestamp 1667941163
transform 1 0 39100 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_421
timestamp 1667941163
transform 1 0 39836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_427
timestamp 1667941163
transform 1 0 40388 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_435
timestamp 1667941163
transform 1 0 41124 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1667941163
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1667941163
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1667941163
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_473
timestamp 1667941163
transform 1 0 44620 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_502
timestamp 1667941163
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1667941163
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1667941163
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_14
timestamp 1667941163
transform 1 0 2392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1667941163
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1667941163
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_261
timestamp 1667941163
transform 1 0 25116 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_268
timestamp 1667941163
transform 1 0 25760 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_280
timestamp 1667941163
transform 1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_291
timestamp 1667941163
transform 1 0 27876 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1667941163
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_317
timestamp 1667941163
transform 1 0 30268 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_337
timestamp 1667941163
transform 1 0 32108 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1667941163
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_371
timestamp 1667941163
transform 1 0 35236 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_379
timestamp 1667941163
transform 1 0 35972 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_400
timestamp 1667941163
transform 1 0 37904 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_414
timestamp 1667941163
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1667941163
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1667941163
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_451
timestamp 1667941163
transform 1 0 42596 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_457
timestamp 1667941163
transform 1 0 43148 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_474
timestamp 1667941163
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_477
timestamp 1667941163
transform 1 0 44988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_485
timestamp 1667941163
transform 1 0 45724 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1667941163
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1667941163
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_513
timestamp 1667941163
transform 1 0 48300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1667941163
transform 1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_16
timestamp 1667941163
transform 1 0 2576 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_28
timestamp 1667941163
transform 1 0 3680 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_40
timestamp 1667941163
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1667941163
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_234
timestamp 1667941163
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_246
timestamp 1667941163
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_258
timestamp 1667941163
transform 1 0 24840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1667941163
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1667941163
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_295
timestamp 1667941163
transform 1 0 28244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_307
timestamp 1667941163
transform 1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_311
timestamp 1667941163
transform 1 0 29716 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_318
timestamp 1667941163
transform 1 0 30360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1667941163
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_367
timestamp 1667941163
transform 1 0 34868 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_377
timestamp 1667941163
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1667941163
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_422
timestamp 1667941163
transform 1 0 39928 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_430
timestamp 1667941163
transform 1 0 40664 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_436
timestamp 1667941163
transform 1 0 41216 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1667941163
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_449
timestamp 1667941163
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_467
timestamp 1667941163
transform 1 0 44068 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_479
timestamp 1667941163
transform 1 0 45172 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_493
timestamp 1667941163
transform 1 0 46460 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_502
timestamp 1667941163
transform 1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_505
timestamp 1667941163
transform 1 0 47564 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_510
timestamp 1667941163
transform 1 0 48024 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1667941163
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_238
timestamp 1667941163
transform 1 0 23000 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_258
timestamp 1667941163
transform 1 0 24840 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_270
timestamp 1667941163
transform 1 0 25944 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_282
timestamp 1667941163
transform 1 0 27048 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_294
timestamp 1667941163
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_327
timestamp 1667941163
transform 1 0 31188 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_335
timestamp 1667941163
transform 1 0 31924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_347
timestamp 1667941163
transform 1 0 33028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_359
timestamp 1667941163
transform 1 0 34132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_379
timestamp 1667941163
transform 1 0 35972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_386
timestamp 1667941163
transform 1 0 36616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_393
timestamp 1667941163
transform 1 0 37260 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_400
timestamp 1667941163
transform 1 0 37904 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_408
timestamp 1667941163
transform 1 0 38640 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1667941163
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1667941163
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1667941163
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_433
timestamp 1667941163
transform 1 0 40940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_437
timestamp 1667941163
transform 1 0 41308 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_442
timestamp 1667941163
transform 1 0 41768 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_449
timestamp 1667941163
transform 1 0 42412 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_461
timestamp 1667941163
transform 1 0 43516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_473
timestamp 1667941163
transform 1 0 44620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_477
timestamp 1667941163
transform 1 0 44988 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_485
timestamp 1667941163
transform 1 0 45724 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_508
timestamp 1667941163
transform 1 0 47840 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_14
timestamp 1667941163
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_26
timestamp 1667941163
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_38
timestamp 1667941163
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1667941163
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_235
timestamp 1667941163
transform 1 0 22724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_247
timestamp 1667941163
transform 1 0 23828 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_265
timestamp 1667941163
transform 1 0 25484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1667941163
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_292
timestamp 1667941163
transform 1 0 27968 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1667941163
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_319
timestamp 1667941163
transform 1 0 30452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_326
timestamp 1667941163
transform 1 0 31096 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1667941163
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_345
timestamp 1667941163
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_357
timestamp 1667941163
transform 1 0 33948 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_369
timestamp 1667941163
transform 1 0 35052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_377
timestamp 1667941163
transform 1 0 35788 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1667941163
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_398
timestamp 1667941163
transform 1 0 37720 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_402
timestamp 1667941163
transform 1 0 38088 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_409
timestamp 1667941163
transform 1 0 38732 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1667941163
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1667941163
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1667941163
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_449
timestamp 1667941163
transform 1 0 42412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_457
timestamp 1667941163
transform 1 0 43148 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_474
timestamp 1667941163
transform 1 0 44712 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_480
timestamp 1667941163
transform 1 0 45264 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_502
timestamp 1667941163
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_505
timestamp 1667941163
transform 1 0 47564 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_510
timestamp 1667941163
transform 1 0 48024 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_273
timestamp 1667941163
transform 1 0 26220 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_279
timestamp 1667941163
transform 1 0 26772 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_291
timestamp 1667941163
transform 1 0 27876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_303
timestamp 1667941163
transform 1 0 28980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_347
timestamp 1667941163
transform 1 0 33028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_351
timestamp 1667941163
transform 1 0 33396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1667941163
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_369
timestamp 1667941163
transform 1 0 35052 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_383
timestamp 1667941163
transform 1 0 36340 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_404
timestamp 1667941163
transform 1 0 38272 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_412
timestamp 1667941163
transform 1 0 39008 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1667941163
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1667941163
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_429
timestamp 1667941163
transform 1 0 40572 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_441
timestamp 1667941163
transform 1 0 41676 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_453
timestamp 1667941163
transform 1 0 42780 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_459
timestamp 1667941163
transform 1 0 43332 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_466
timestamp 1667941163
transform 1 0 43976 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_474
timestamp 1667941163
transform 1 0 44712 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1667941163
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_489
timestamp 1667941163
transform 1 0 46092 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_514
timestamp 1667941163
transform 1 0 48392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_244
timestamp 1667941163
transform 1 0 23552 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_256
timestamp 1667941163
transform 1 0 24656 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1667941163
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1667941163
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_291
timestamp 1667941163
transform 1 0 27876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_303
timestamp 1667941163
transform 1 0 28980 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_311
timestamp 1667941163
transform 1 0 29716 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_326
timestamp 1667941163
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1667941163
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_345
timestamp 1667941163
transform 1 0 32844 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_362
timestamp 1667941163
transform 1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_370
timestamp 1667941163
transform 1 0 35144 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1667941163
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1667941163
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1667941163
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1667941163
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1667941163
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_449
timestamp 1667941163
transform 1 0 42412 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_457
timestamp 1667941163
transform 1 0 43148 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_463
timestamp 1667941163
transform 1 0 43700 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_475
timestamp 1667941163
transform 1 0 44804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_483
timestamp 1667941163
transform 1 0 45540 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_502
timestamp 1667941163
transform 1 0 47288 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_505
timestamp 1667941163
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_510
timestamp 1667941163
transform 1 0 48024 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1667941163
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1667941163
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1667941163
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1667941163
transform 1 0 27048 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_296
timestamp 1667941163
transform 1 0 28336 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_329
timestamp 1667941163
transform 1 0 31372 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_338
timestamp 1667941163
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_350
timestamp 1667941163
transform 1 0 33304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1667941163
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_373
timestamp 1667941163
transform 1 0 35420 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_385
timestamp 1667941163
transform 1 0 36524 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_397
timestamp 1667941163
transform 1 0 37628 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_409
timestamp 1667941163
transform 1 0 38732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1667941163
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_421
timestamp 1667941163
transform 1 0 39836 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_428
timestamp 1667941163
transform 1 0 40480 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_440
timestamp 1667941163
transform 1 0 41584 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_446
timestamp 1667941163
transform 1 0 42136 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_454
timestamp 1667941163
transform 1 0 42872 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_459
timestamp 1667941163
transform 1 0 43332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_468
timestamp 1667941163
transform 1 0 44160 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_477
timestamp 1667941163
transform 1 0 44988 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_490
timestamp 1667941163
transform 1 0 46184 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_498
timestamp 1667941163
transform 1 0 46920 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_510
timestamp 1667941163
transform 1 0 48024 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_233
timestamp 1667941163
transform 1 0 22540 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_241
timestamp 1667941163
transform 1 0 23276 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_254
timestamp 1667941163
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_263
timestamp 1667941163
transform 1 0 25300 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_271
timestamp 1667941163
transform 1 0 26036 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1667941163
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_302
timestamp 1667941163
transform 1 0 28888 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_314
timestamp 1667941163
transform 1 0 29992 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_322
timestamp 1667941163
transform 1 0 30728 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_328
timestamp 1667941163
transform 1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_343
timestamp 1667941163
transform 1 0 32660 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_350
timestamp 1667941163
transform 1 0 33304 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_362
timestamp 1667941163
transform 1 0 34408 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_376
timestamp 1667941163
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1667941163
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_399
timestamp 1667941163
transform 1 0 37812 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1667941163
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_423
timestamp 1667941163
transform 1 0 40020 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_429
timestamp 1667941163
transform 1 0 40572 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1667941163
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_449
timestamp 1667941163
transform 1 0 42412 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_453
timestamp 1667941163
transform 1 0 42780 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_470
timestamp 1667941163
transform 1 0 44344 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_482
timestamp 1667941163
transform 1 0 45448 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_488
timestamp 1667941163
transform 1 0 46000 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_495
timestamp 1667941163
transform 1 0 46644 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1667941163
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_505
timestamp 1667941163
transform 1 0 47564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_510
timestamp 1667941163
transform 1 0 48024 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_237
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1667941163
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_260
timestamp 1667941163
transform 1 0 25024 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_268
timestamp 1667941163
transform 1 0 25760 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_274
timestamp 1667941163
transform 1 0 26312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_285
timestamp 1667941163
transform 1 0 27324 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_292
timestamp 1667941163
transform 1 0 27968 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1667941163
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_315
timestamp 1667941163
transform 1 0 30084 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_343
timestamp 1667941163
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 1667941163
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_369
timestamp 1667941163
transform 1 0 35052 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_379
timestamp 1667941163
transform 1 0 35972 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1667941163
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1667941163
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_421
timestamp 1667941163
transform 1 0 39836 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_427
timestamp 1667941163
transform 1 0 40388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_443
timestamp 1667941163
transform 1 0 41860 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_450
timestamp 1667941163
transform 1 0 42504 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_462
timestamp 1667941163
transform 1 0 43608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1667941163
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1667941163
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_477
timestamp 1667941163
transform 1 0 44988 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_489
timestamp 1667941163
transform 1 0 46092 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_514
timestamp 1667941163
transform 1 0 48392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_256
timestamp 1667941163
transform 1 0 24656 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_268
timestamp 1667941163
transform 1 0 25760 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_274
timestamp 1667941163
transform 1 0 26312 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1667941163
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_291
timestamp 1667941163
transform 1 0 27876 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_299
timestamp 1667941163
transform 1 0 28612 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_316
timestamp 1667941163
transform 1 0 30176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_326
timestamp 1667941163
transform 1 0 31096 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1667941163
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_357
timestamp 1667941163
transform 1 0 33948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_366
timestamp 1667941163
transform 1 0 34776 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_377
timestamp 1667941163
transform 1 0 35788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_387
timestamp 1667941163
transform 1 0 36708 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_411
timestamp 1667941163
transform 1 0 38916 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_426
timestamp 1667941163
transform 1 0 40296 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_433
timestamp 1667941163
transform 1 0 40940 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_441
timestamp 1667941163
transform 1 0 41676 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_446
timestamp 1667941163
transform 1 0 42136 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_449
timestamp 1667941163
transform 1 0 42412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_453
timestamp 1667941163
transform 1 0 42780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_460
timestamp 1667941163
transform 1 0 43424 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_467
timestamp 1667941163
transform 1 0 44068 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_479
timestamp 1667941163
transform 1 0 45172 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_499
timestamp 1667941163
transform 1 0 47012 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1667941163
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_505
timestamp 1667941163
transform 1 0 47564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_510
timestamp 1667941163
transform 1 0 48024 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_238
timestamp 1667941163
transform 1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1667941163
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_271
timestamp 1667941163
transform 1 0 26036 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_278
timestamp 1667941163
transform 1 0 26680 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1667941163
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_327
timestamp 1667941163
transform 1 0 31188 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_344
timestamp 1667941163
transform 1 0 32752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1667941163
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_375
timestamp 1667941163
transform 1 0 35604 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_384
timestamp 1667941163
transform 1 0 36432 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_396
timestamp 1667941163
transform 1 0 37536 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_408
timestamp 1667941163
transform 1 0 38640 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1667941163
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_421
timestamp 1667941163
transform 1 0 39836 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_430
timestamp 1667941163
transform 1 0 40664 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_442
timestamp 1667941163
transform 1 0 41768 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_457
timestamp 1667941163
transform 1 0 43148 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_468
timestamp 1667941163
transform 1 0 44160 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_477
timestamp 1667941163
transform 1 0 44988 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_483
timestamp 1667941163
transform 1 0 45540 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_487
timestamp 1667941163
transform 1 0 45908 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_514
timestamp 1667941163
transform 1 0 48392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_265
timestamp 1667941163
transform 1 0 25484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1667941163
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1667941163
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_344
timestamp 1667941163
transform 1 0 32752 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_351
timestamp 1667941163
transform 1 0 33396 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_363
timestamp 1667941163
transform 1 0 34500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_371
timestamp 1667941163
transform 1 0 35236 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_375
timestamp 1667941163
transform 1 0 35604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_387
timestamp 1667941163
transform 1 0 36708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_409
timestamp 1667941163
transform 1 0 38732 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_414
timestamp 1667941163
transform 1 0 39192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_425
timestamp 1667941163
transform 1 0 40204 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_436
timestamp 1667941163
transform 1 0 41216 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_449
timestamp 1667941163
transform 1 0 42412 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_471
timestamp 1667941163
transform 1 0 44436 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_484
timestamp 1667941163
transform 1 0 45632 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_494
timestamp 1667941163
transform 1 0 46552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_498
timestamp 1667941163
transform 1 0 46920 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_502
timestamp 1667941163
transform 1 0 47288 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_505
timestamp 1667941163
transform 1 0 47564 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_510
timestamp 1667941163
transform 1 0 48024 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_273
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_281
timestamp 1667941163
transform 1 0 26956 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_293
timestamp 1667941163
transform 1 0 28060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1667941163
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_316
timestamp 1667941163
transform 1 0 30176 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_324
timestamp 1667941163
transform 1 0 30912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_332
timestamp 1667941163
transform 1 0 31648 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_354
timestamp 1667941163
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1667941163
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_383
timestamp 1667941163
transform 1 0 36340 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_411
timestamp 1667941163
transform 1 0 38916 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1667941163
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_421
timestamp 1667941163
transform 1 0 39836 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_425
timestamp 1667941163
transform 1 0 40204 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_432
timestamp 1667941163
transform 1 0 40848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_444
timestamp 1667941163
transform 1 0 41952 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_452
timestamp 1667941163
transform 1 0 42688 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_462
timestamp 1667941163
transform 1 0 43608 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_474
timestamp 1667941163
transform 1 0 44712 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_477
timestamp 1667941163
transform 1 0 44988 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_487
timestamp 1667941163
transform 1 0 45908 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_494
timestamp 1667941163
transform 1 0 46552 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_506
timestamp 1667941163
transform 1 0 47656 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_514
timestamp 1667941163
transform 1 0 48392 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_254
timestamp 1667941163
transform 1 0 24472 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_269
timestamp 1667941163
transform 1 0 25852 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_292
timestamp 1667941163
transform 1 0 27968 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_303
timestamp 1667941163
transform 1 0 28980 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_323
timestamp 1667941163
transform 1 0 30820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_327
timestamp 1667941163
transform 1 0 31188 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1667941163
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_346
timestamp 1667941163
transform 1 0 32936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_374
timestamp 1667941163
transform 1 0 35512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_381
timestamp 1667941163
transform 1 0 36156 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1667941163
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_398
timestamp 1667941163
transform 1 0 37720 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_410
timestamp 1667941163
transform 1 0 38824 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_422
timestamp 1667941163
transform 1 0 39928 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_430
timestamp 1667941163
transform 1 0 40664 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_437
timestamp 1667941163
transform 1 0 41308 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_445
timestamp 1667941163
transform 1 0 42044 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1667941163
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1667941163
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1667941163
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1667941163
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_501
timestamp 1667941163
transform 1 0 47196 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1667941163
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1667941163
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_271
timestamp 1667941163
transform 1 0 26036 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_278
timestamp 1667941163
transform 1 0 26680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_285
timestamp 1667941163
transform 1 0 27324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1667941163
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_315
timestamp 1667941163
transform 1 0 30084 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_372
timestamp 1667941163
transform 1 0 35328 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_400
timestamp 1667941163
transform 1 0 37904 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_410
timestamp 1667941163
transform 1 0 38824 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_414
timestamp 1667941163
transform 1 0 39192 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1667941163
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_421
timestamp 1667941163
transform 1 0 39836 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_428
timestamp 1667941163
transform 1 0 40480 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_439
timestamp 1667941163
transform 1 0 41492 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_451
timestamp 1667941163
transform 1 0 42596 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_463
timestamp 1667941163
transform 1 0 43700 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_470
timestamp 1667941163
transform 1 0 44344 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_477
timestamp 1667941163
transform 1 0 44988 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_485
timestamp 1667941163
transform 1 0 45724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_497
timestamp 1667941163
transform 1 0 46828 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_514
timestamp 1667941163
transform 1 0 48392 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_11
timestamp 1667941163
transform 1 0 2116 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_16
timestamp 1667941163
transform 1 0 2576 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_28
timestamp 1667941163
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_40
timestamp 1667941163
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1667941163
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_266
timestamp 1667941163
transform 1 0 25576 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1667941163
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_289
timestamp 1667941163
transform 1 0 27692 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_297
timestamp 1667941163
transform 1 0 28428 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_316
timestamp 1667941163
transform 1 0 30176 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_328
timestamp 1667941163
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_347
timestamp 1667941163
transform 1 0 33028 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_359
timestamp 1667941163
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_371
timestamp 1667941163
transform 1 0 35236 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_383
timestamp 1667941163
transform 1 0 36340 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_399
timestamp 1667941163
transform 1 0 37812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_407
timestamp 1667941163
transform 1 0 38548 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_416
timestamp 1667941163
transform 1 0 39376 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_429
timestamp 1667941163
transform 1 0 40572 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_442
timestamp 1667941163
transform 1 0 41768 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_449
timestamp 1667941163
transform 1 0 42412 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_454
timestamp 1667941163
transform 1 0 42872 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_466
timestamp 1667941163
transform 1 0 43976 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_474
timestamp 1667941163
transform 1 0 44712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_483
timestamp 1667941163
transform 1 0 45540 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_494
timestamp 1667941163
transform 1 0 46552 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_502
timestamp 1667941163
transform 1 0 47288 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_505
timestamp 1667941163
transform 1 0 47564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_510
timestamp 1667941163
transform 1 0 48024 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1667941163
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_271
timestamp 1667941163
transform 1 0 26036 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_281
timestamp 1667941163
transform 1 0 26956 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_293
timestamp 1667941163
transform 1 0 28060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1667941163
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_314
timestamp 1667941163
transform 1 0 29992 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_326
timestamp 1667941163
transform 1 0 31096 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_353
timestamp 1667941163
transform 1 0 33580 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1667941163
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_399
timestamp 1667941163
transform 1 0 37812 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_417
timestamp 1667941163
transform 1 0 39468 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_421
timestamp 1667941163
transform 1 0 39836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_434
timestamp 1667941163
transform 1 0 41032 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_438
timestamp 1667941163
transform 1 0 41400 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_455
timestamp 1667941163
transform 1 0 42964 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_466
timestamp 1667941163
transform 1 0 43976 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_473
timestamp 1667941163
transform 1 0 44620 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_477
timestamp 1667941163
transform 1 0 44988 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_486
timestamp 1667941163
transform 1 0 45816 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_492
timestamp 1667941163
transform 1 0 46368 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_514
timestamp 1667941163
transform 1 0 48392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_14
timestamp 1667941163
transform 1 0 2392 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_26
timestamp 1667941163
transform 1 0 3496 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_38
timestamp 1667941163
transform 1 0 4600 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_50
timestamp 1667941163
transform 1 0 5704 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_254
timestamp 1667941163
transform 1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_263
timestamp 1667941163
transform 1 0 25300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1667941163
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_286
timestamp 1667941163
transform 1 0 27416 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_298
timestamp 1667941163
transform 1 0 28520 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_310
timestamp 1667941163
transform 1 0 29624 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_322
timestamp 1667941163
transform 1 0 30728 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1667941163
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_356
timestamp 1667941163
transform 1 0 33856 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_376
timestamp 1667941163
transform 1 0 35696 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1667941163
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1667941163
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_410
timestamp 1667941163
transform 1 0 38824 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_422
timestamp 1667941163
transform 1 0 39928 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_430
timestamp 1667941163
transform 1 0 40664 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_435
timestamp 1667941163
transform 1 0 41124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1667941163
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1667941163
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1667941163
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_473
timestamp 1667941163
transform 1 0 44620 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_477
timestamp 1667941163
transform 1 0 44988 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1667941163
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1667941163
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1667941163
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_505
timestamp 1667941163
transform 1 0 47564 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_510
timestamp 1667941163
transform 1 0 48024 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_287
timestamp 1667941163
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_299
timestamp 1667941163
transform 1 0 28612 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1667941163
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_316
timestamp 1667941163
transform 1 0 30176 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_331
timestamp 1667941163
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_343
timestamp 1667941163
transform 1 0 32660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_355
timestamp 1667941163
transform 1 0 33764 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1667941163
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_372
timestamp 1667941163
transform 1 0 35328 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_379
timestamp 1667941163
transform 1 0 35972 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1667941163
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1667941163
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1667941163
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_421
timestamp 1667941163
transform 1 0 39836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_426
timestamp 1667941163
transform 1 0 40296 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1667941163
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1667941163
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_457
timestamp 1667941163
transform 1 0 43148 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_465
timestamp 1667941163
transform 1 0 43884 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1667941163
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1667941163
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1667941163
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1667941163
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_501
timestamp 1667941163
transform 1 0 47196 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_509
timestamp 1667941163
transform 1 0 47932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_514
timestamp 1667941163
transform 1 0 48392 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_245
timestamp 1667941163
transform 1 0 23644 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_264
timestamp 1667941163
transform 1 0 25392 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1667941163
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_288
timestamp 1667941163
transform 1 0 27600 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_294
timestamp 1667941163
transform 1 0 28152 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_311
timestamp 1667941163
transform 1 0 29716 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1667941163
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_353
timestamp 1667941163
transform 1 0 33580 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_359
timestamp 1667941163
transform 1 0 34132 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_379
timestamp 1667941163
transform 1 0 35972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_401
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_408
timestamp 1667941163
transform 1 0 38640 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_414
timestamp 1667941163
transform 1 0 39192 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_421
timestamp 1667941163
transform 1 0 39836 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_429
timestamp 1667941163
transform 1 0 40572 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_437
timestamp 1667941163
transform 1 0 41308 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_445
timestamp 1667941163
transform 1 0 42044 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_449
timestamp 1667941163
transform 1 0 42412 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_462
timestamp 1667941163
transform 1 0 43608 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_466
timestamp 1667941163
transform 1 0 43976 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_473
timestamp 1667941163
transform 1 0 44620 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_481
timestamp 1667941163
transform 1 0 45356 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_491
timestamp 1667941163
transform 1 0 46276 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_59_501
timestamp 1667941163
transform 1 0 47196 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1667941163
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1667941163
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_282
timestamp 1667941163
transform 1 0 27048 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_294
timestamp 1667941163
transform 1 0 28152 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_302
timestamp 1667941163
transform 1 0 28888 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1667941163
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_316
timestamp 1667941163
transform 1 0 30176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_325
timestamp 1667941163
transform 1 0 31004 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_332
timestamp 1667941163
transform 1 0 31648 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_340
timestamp 1667941163
transform 1 0 32384 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_344
timestamp 1667941163
transform 1 0 32752 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_353
timestamp 1667941163
transform 1 0 33580 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_361
timestamp 1667941163
transform 1 0 34316 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_397
timestamp 1667941163
transform 1 0 37628 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1667941163
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_411
timestamp 1667941163
transform 1 0 38916 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1667941163
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_421
timestamp 1667941163
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_429
timestamp 1667941163
transform 1 0 40572 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_441
timestamp 1667941163
transform 1 0 41676 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_453
timestamp 1667941163
transform 1 0 42780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_462
timestamp 1667941163
transform 1 0 43608 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_473
timestamp 1667941163
transform 1 0 44620 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_477
timestamp 1667941163
transform 1 0 44988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_488
timestamp 1667941163
transform 1 0 46000 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_496
timestamp 1667941163
transform 1 0 46736 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_514
timestamp 1667941163
transform 1 0 48392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_271
timestamp 1667941163
transform 1 0 26036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_288
timestamp 1667941163
transform 1 0 27600 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_300
timestamp 1667941163
transform 1 0 28704 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_304
timestamp 1667941163
transform 1 0 29072 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_321
timestamp 1667941163
transform 1 0 30636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1667941163
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_355
timestamp 1667941163
transform 1 0 33764 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_368
timestamp 1667941163
transform 1 0 34960 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_376
timestamp 1667941163
transform 1 0 35696 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_381
timestamp 1667941163
transform 1 0 36156 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1667941163
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_401
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_411
timestamp 1667941163
transform 1 0 38916 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_424
timestamp 1667941163
transform 1 0 40112 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_435
timestamp 1667941163
transform 1 0 41124 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_444
timestamp 1667941163
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_449
timestamp 1667941163
transform 1 0 42412 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_469
timestamp 1667941163
transform 1 0 44252 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_478
timestamp 1667941163
transform 1 0 45080 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_490
timestamp 1667941163
transform 1 0 46184 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_494
timestamp 1667941163
transform 1 0 46552 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_499
timestamp 1667941163
transform 1 0 47012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1667941163
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1667941163
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1667941163
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_239
timestamp 1667941163
transform 1 0 23092 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_243
timestamp 1667941163
transform 1 0 23460 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1667941163
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_291
timestamp 1667941163
transform 1 0 27876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1667941163
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1667941163
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_347
timestamp 1667941163
transform 1 0 33028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_359
timestamp 1667941163
transform 1 0 34132 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_409
timestamp 1667941163
transform 1 0 38732 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_416
timestamp 1667941163
transform 1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_421
timestamp 1667941163
transform 1 0 39836 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_429
timestamp 1667941163
transform 1 0 40572 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_436
timestamp 1667941163
transform 1 0 41216 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_460
timestamp 1667941163
transform 1 0 43424 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_466
timestamp 1667941163
transform 1 0 43976 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_470
timestamp 1667941163
transform 1 0 44344 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1667941163
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_489
timestamp 1667941163
transform 1 0 46092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_514
timestamp 1667941163
transform 1 0 48392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_255
timestamp 1667941163
transform 1 0 24564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_264
timestamp 1667941163
transform 1 0 25392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1667941163
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_299
timestamp 1667941163
transform 1 0 28612 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_311
timestamp 1667941163
transform 1 0 29716 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_321
timestamp 1667941163
transform 1 0 30636 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1667941163
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_345
timestamp 1667941163
transform 1 0 32844 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_354
timestamp 1667941163
transform 1 0 33672 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_360
timestamp 1667941163
transform 1 0 34224 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_377
timestamp 1667941163
transform 1 0 35788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1667941163
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_400
timestamp 1667941163
transform 1 0 37904 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_432
timestamp 1667941163
transform 1 0 40848 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1667941163
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1667941163
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_449
timestamp 1667941163
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_454
timestamp 1667941163
transform 1 0 42872 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_466
timestamp 1667941163
transform 1 0 43976 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_478
timestamp 1667941163
transform 1 0 45080 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_490
timestamp 1667941163
transform 1 0 46184 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_498
timestamp 1667941163
transform 1 0 46920 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_502
timestamp 1667941163
transform 1 0 47288 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_505
timestamp 1667941163
transform 1 0 47564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_510
timestamp 1667941163
transform 1 0 48024 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1667941163
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1667941163
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1667941163
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1667941163
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1667941163
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_260
timestamp 1667941163
transform 1 0 25024 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_268
timestamp 1667941163
transform 1 0 25760 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_276
timestamp 1667941163
transform 1 0 26496 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_288
timestamp 1667941163
transform 1 0 27600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_297
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1667941163
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_333
timestamp 1667941163
transform 1 0 31740 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_340
timestamp 1667941163
transform 1 0 32384 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_346
timestamp 1667941163
transform 1 0 32936 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_354
timestamp 1667941163
transform 1 0 33672 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_375
timestamp 1667941163
transform 1 0 35604 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_384
timestamp 1667941163
transform 1 0 36432 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_396
timestamp 1667941163
transform 1 0 37536 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_404
timestamp 1667941163
transform 1 0 38272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_416
timestamp 1667941163
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1667941163
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_431
timestamp 1667941163
transform 1 0 40756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_441
timestamp 1667941163
transform 1 0 41676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_461
timestamp 1667941163
transform 1 0 43516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_470
timestamp 1667941163
transform 1 0 44344 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_477
timestamp 1667941163
transform 1 0 44988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_481
timestamp 1667941163
transform 1 0 45356 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_487
timestamp 1667941163
transform 1 0 45908 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_514
timestamp 1667941163
transform 1 0 48392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1667941163
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1667941163
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1667941163
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1667941163
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1667941163
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1667941163
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1667941163
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1667941163
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1667941163
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1667941163
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1667941163
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1667941163
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1667941163
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1667941163
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1667941163
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1667941163
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1667941163
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1667941163
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1667941163
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1667941163
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1667941163
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1667941163
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1667941163
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1667941163
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1667941163
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_237
timestamp 1667941163
transform 1 0 22908 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_243
timestamp 1667941163
transform 1 0 23460 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_260
timestamp 1667941163
transform 1 0 25024 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_272
timestamp 1667941163
transform 1 0 26128 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1667941163
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_309
timestamp 1667941163
transform 1 0 29532 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_321
timestamp 1667941163
transform 1 0 30636 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_330
timestamp 1667941163
transform 1 0 31464 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_337
timestamp 1667941163
transform 1 0 32108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_341
timestamp 1667941163
transform 1 0 32476 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_358
timestamp 1667941163
transform 1 0 34040 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_370
timestamp 1667941163
transform 1 0 35144 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_382
timestamp 1667941163
transform 1 0 36248 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_386
timestamp 1667941163
transform 1 0 36616 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_390
timestamp 1667941163
transform 1 0 36984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 1667941163
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_411
timestamp 1667941163
transform 1 0 38916 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_435
timestamp 1667941163
transform 1 0 41124 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1667941163
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_449
timestamp 1667941163
transform 1 0 42412 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_455
timestamp 1667941163
transform 1 0 42964 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_459
timestamp 1667941163
transform 1 0 43332 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_479
timestamp 1667941163
transform 1 0 45172 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_487
timestamp 1667941163
transform 1 0 45908 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_492
timestamp 1667941163
transform 1 0 46368 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_499
timestamp 1667941163
transform 1 0 47012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1667941163
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_505
timestamp 1667941163
transform 1 0 47564 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_510
timestamp 1667941163
transform 1 0 48024 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1667941163
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1667941163
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1667941163
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1667941163
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1667941163
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1667941163
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1667941163
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1667941163
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1667941163
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1667941163
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1667941163
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1667941163
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1667941163
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1667941163
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1667941163
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1667941163
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1667941163
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1667941163
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1667941163
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1667941163
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1667941163
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1667941163
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1667941163
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1667941163
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1667941163
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1667941163
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1667941163
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1667941163
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_258
timestamp 1667941163
transform 1 0 24840 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_264
timestamp 1667941163
transform 1 0 25392 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_271
timestamp 1667941163
transform 1 0 26036 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_283
timestamp 1667941163
transform 1 0 27140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_295
timestamp 1667941163
transform 1 0 28244 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1667941163
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1667941163
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1667941163
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_321
timestamp 1667941163
transform 1 0 30636 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_339
timestamp 1667941163
transform 1 0 32292 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_348
timestamp 1667941163
transform 1 0 33120 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_355
timestamp 1667941163
transform 1 0 33764 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1667941163
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1667941163
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1667941163
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_394
timestamp 1667941163
transform 1 0 37352 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_406
timestamp 1667941163
transform 1 0 38456 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_415
timestamp 1667941163
transform 1 0 39284 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1667941163
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_421
timestamp 1667941163
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_426
timestamp 1667941163
transform 1 0 40296 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_446
timestamp 1667941163
transform 1 0 42136 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_458
timestamp 1667941163
transform 1 0 43240 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_466
timestamp 1667941163
transform 1 0 43976 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_474
timestamp 1667941163
transform 1 0 44712 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_477
timestamp 1667941163
transform 1 0 44988 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_484
timestamp 1667941163
transform 1 0 45632 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_492
timestamp 1667941163
transform 1 0 46368 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_514
timestamp 1667941163
transform 1 0 48392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1667941163
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1667941163
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1667941163
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1667941163
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1667941163
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1667941163
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1667941163
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1667941163
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1667941163
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1667941163
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1667941163
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1667941163
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1667941163
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1667941163
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1667941163
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1667941163
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1667941163
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1667941163
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1667941163
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1667941163
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1667941163
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1667941163
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1667941163
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1667941163
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1667941163
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1667941163
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1667941163
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_261
timestamp 1667941163
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_271
timestamp 1667941163
transform 1 0 26036 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1667941163
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1667941163
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_309
timestamp 1667941163
transform 1 0 29532 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_321
timestamp 1667941163
transform 1 0 30636 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_328
timestamp 1667941163
transform 1 0 31280 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_337
timestamp 1667941163
transform 1 0 32108 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_343
timestamp 1667941163
transform 1 0 32660 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_351
timestamp 1667941163
transform 1 0 33396 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_363
timestamp 1667941163
transform 1 0 34500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_371
timestamp 1667941163
transform 1 0 35236 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_389
timestamp 1667941163
transform 1 0 36892 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_393
timestamp 1667941163
transform 1 0 37260 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_397
timestamp 1667941163
transform 1 0 37628 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_404
timestamp 1667941163
transform 1 0 38272 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_412
timestamp 1667941163
transform 1 0 39008 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1667941163
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1667941163
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1667941163
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1667941163
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_449
timestamp 1667941163
transform 1 0 42412 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_457
timestamp 1667941163
transform 1 0 43148 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_464
timestamp 1667941163
transform 1 0 43792 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_474
timestamp 1667941163
transform 1 0 44712 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_478
timestamp 1667941163
transform 1 0 45080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_482
timestamp 1667941163
transform 1 0 45448 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_502
timestamp 1667941163
transform 1 0 47288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_505
timestamp 1667941163
transform 1 0 47564 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_510
timestamp 1667941163
transform 1 0 48024 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1667941163
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1667941163
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1667941163
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1667941163
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1667941163
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1667941163
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1667941163
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1667941163
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1667941163
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1667941163
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1667941163
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1667941163
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1667941163
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1667941163
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1667941163
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1667941163
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1667941163
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1667941163
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1667941163
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1667941163
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1667941163
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1667941163
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1667941163
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1667941163
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1667941163
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_245
timestamp 1667941163
transform 1 0 23644 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1667941163
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1667941163
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_260
timestamp 1667941163
transform 1 0 25024 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_264
timestamp 1667941163
transform 1 0 25392 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_281
timestamp 1667941163
transform 1 0 26956 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_285
timestamp 1667941163
transform 1 0 27324 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_291
timestamp 1667941163
transform 1 0 27876 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_303
timestamp 1667941163
transform 1 0 28980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1667941163
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1667941163
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_316
timestamp 1667941163
transform 1 0 30176 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_328
timestamp 1667941163
transform 1 0 31280 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_334
timestamp 1667941163
transform 1 0 31832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_340
timestamp 1667941163
transform 1 0 32384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_344
timestamp 1667941163
transform 1 0 32752 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_348
timestamp 1667941163
transform 1 0 33120 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1667941163
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_365
timestamp 1667941163
transform 1 0 34684 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_374
timestamp 1667941163
transform 1 0 35512 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_390
timestamp 1667941163
transform 1 0 36984 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_418
timestamp 1667941163
transform 1 0 39560 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1667941163
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1667941163
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_445
timestamp 1667941163
transform 1 0 42044 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_451
timestamp 1667941163
transform 1 0 42596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_463
timestamp 1667941163
transform 1 0 43700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1667941163
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_477
timestamp 1667941163
transform 1 0 44988 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_482
timestamp 1667941163
transform 1 0 45448 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_490
timestamp 1667941163
transform 1 0 46184 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_514
timestamp 1667941163
transform 1 0 48392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1667941163
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1667941163
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1667941163
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1667941163
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1667941163
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1667941163
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1667941163
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1667941163
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1667941163
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1667941163
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1667941163
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1667941163
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1667941163
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1667941163
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1667941163
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1667941163
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1667941163
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1667941163
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1667941163
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1667941163
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1667941163
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1667941163
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1667941163
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1667941163
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1667941163
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_237
timestamp 1667941163
transform 1 0 22908 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_261
timestamp 1667941163
transform 1 0 25116 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_265
timestamp 1667941163
transform 1 0 25484 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_271
timestamp 1667941163
transform 1 0 26036 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1667941163
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_281
timestamp 1667941163
transform 1 0 26956 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_289
timestamp 1667941163
transform 1 0 27692 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_295
timestamp 1667941163
transform 1 0 28244 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_315
timestamp 1667941163
transform 1 0 30084 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_326
timestamp 1667941163
transform 1 0 31096 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 1667941163
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_337
timestamp 1667941163
transform 1 0 32108 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_345
timestamp 1667941163
transform 1 0 32844 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_364
timestamp 1667941163
transform 1 0 34592 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_378
timestamp 1667941163
transform 1 0 35880 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_389
timestamp 1667941163
transform 1 0 36892 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1667941163
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_405
timestamp 1667941163
transform 1 0 38364 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_424
timestamp 1667941163
transform 1 0 40112 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_436
timestamp 1667941163
transform 1 0 41216 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_443
timestamp 1667941163
transform 1 0 41860 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1667941163
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_449
timestamp 1667941163
transform 1 0 42412 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_458
timestamp 1667941163
transform 1 0 43240 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_464
timestamp 1667941163
transform 1 0 43792 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_470
timestamp 1667941163
transform 1 0 44344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_490
timestamp 1667941163
transform 1 0 46184 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_498
timestamp 1667941163
transform 1 0 46920 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_502
timestamp 1667941163
transform 1 0 47288 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_505
timestamp 1667941163
transform 1 0 47564 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_510
timestamp 1667941163
transform 1 0 48024 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_3
timestamp 1667941163
transform 1 0 1380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_11
timestamp 1667941163
transform 1 0 2116 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_16
timestamp 1667941163
transform 1 0 2576 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1667941163
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1667941163
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1667941163
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1667941163
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1667941163
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1667941163
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1667941163
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1667941163
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1667941163
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1667941163
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1667941163
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1667941163
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1667941163
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1667941163
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1667941163
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1667941163
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1667941163
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1667941163
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1667941163
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1667941163
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1667941163
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1667941163
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_245
timestamp 1667941163
transform 1 0 23644 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1667941163
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1667941163
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_260
timestamp 1667941163
transform 1 0 25024 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_272
timestamp 1667941163
transform 1 0 26128 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_284
timestamp 1667941163
transform 1 0 27232 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_296
timestamp 1667941163
transform 1 0 28336 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_303
timestamp 1667941163
transform 1 0 28980 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1667941163
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1667941163
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_316
timestamp 1667941163
transform 1 0 30176 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_328
timestamp 1667941163
transform 1 0 31280 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_340
timestamp 1667941163
transform 1 0 32384 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_362
timestamp 1667941163
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_365
timestamp 1667941163
transform 1 0 34684 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_373
timestamp 1667941163
transform 1 0 35420 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_379
timestamp 1667941163
transform 1 0 35972 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_387
timestamp 1667941163
transform 1 0 36708 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_396
timestamp 1667941163
transform 1 0 37536 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_408
timestamp 1667941163
transform 1 0 38640 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_70_417
timestamp 1667941163
transform 1 0 39468 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_421
timestamp 1667941163
transform 1 0 39836 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_428
timestamp 1667941163
transform 1 0 40480 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_448
timestamp 1667941163
transform 1 0 42320 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_468
timestamp 1667941163
transform 1 0 44160 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_477
timestamp 1667941163
transform 1 0 44988 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_484
timestamp 1667941163
transform 1 0 45632 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_492
timestamp 1667941163
transform 1 0 46368 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_514
timestamp 1667941163
transform 1 0 48392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1667941163
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1667941163
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_31
timestamp 1667941163
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_43
timestamp 1667941163
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1667941163
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1667941163
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1667941163
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1667941163
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1667941163
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1667941163
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1667941163
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1667941163
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1667941163
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1667941163
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1667941163
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1667941163
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1667941163
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1667941163
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1667941163
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1667941163
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1667941163
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1667941163
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1667941163
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1667941163
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1667941163
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_249
timestamp 1667941163
transform 1 0 24012 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_267
timestamp 1667941163
transform 1 0 25668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1667941163
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1667941163
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1667941163
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1667941163
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_317
timestamp 1667941163
transform 1 0 30268 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_326
timestamp 1667941163
transform 1 0 31096 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_334
timestamp 1667941163
transform 1 0 31832 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_337
timestamp 1667941163
transform 1 0 32108 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_344
timestamp 1667941163
transform 1 0 32752 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_352
timestamp 1667941163
transform 1 0 33488 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_358
timestamp 1667941163
transform 1 0 34040 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_370
timestamp 1667941163
transform 1 0 35144 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_382
timestamp 1667941163
transform 1 0 36248 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_390
timestamp 1667941163
transform 1 0 36984 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_393
timestamp 1667941163
transform 1 0 37260 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_401
timestamp 1667941163
transform 1 0 37996 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_419
timestamp 1667941163
transform 1 0 39652 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_426
timestamp 1667941163
transform 1 0 40296 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_437
timestamp 1667941163
transform 1 0 41308 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_446
timestamp 1667941163
transform 1 0 42136 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_449
timestamp 1667941163
transform 1 0 42412 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_459
timestamp 1667941163
transform 1 0 43332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_471
timestamp 1667941163
transform 1 0 44436 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_489
timestamp 1667941163
transform 1 0 46092 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_497
timestamp 1667941163
transform 1 0 46828 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_502
timestamp 1667941163
transform 1 0 47288 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_505
timestamp 1667941163
transform 1 0 47564 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_510
timestamp 1667941163
transform 1 0 48024 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_72_3
timestamp 1667941163
transform 1 0 1380 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_14
timestamp 1667941163
transform 1 0 2392 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1667941163
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1667941163
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1667941163
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1667941163
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1667941163
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1667941163
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1667941163
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1667941163
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1667941163
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1667941163
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1667941163
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1667941163
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1667941163
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1667941163
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1667941163
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1667941163
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1667941163
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1667941163
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1667941163
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1667941163
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1667941163
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1667941163
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1667941163
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1667941163
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1667941163
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1667941163
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_271
timestamp 1667941163
transform 1 0 26036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_277
timestamp 1667941163
transform 1 0 26588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_294
timestamp 1667941163
transform 1 0 28152 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_303
timestamp 1667941163
transform 1 0 28980 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1667941163
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_309
timestamp 1667941163
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_317
timestamp 1667941163
transform 1 0 30268 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_327
timestamp 1667941163
transform 1 0 31188 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_347
timestamp 1667941163
transform 1 0 33028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_359
timestamp 1667941163
transform 1 0 34132 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1667941163
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1667941163
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_372
timestamp 1667941163
transform 1 0 35328 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_380
timestamp 1667941163
transform 1 0 36064 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_399
timestamp 1667941163
transform 1 0 37812 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_408
timestamp 1667941163
transform 1 0 38640 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1667941163
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1667941163
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_445
timestamp 1667941163
transform 1 0 42044 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_451
timestamp 1667941163
transform 1 0 42596 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_457
timestamp 1667941163
transform 1 0 43148 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_464
timestamp 1667941163
transform 1 0 43792 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_477
timestamp 1667941163
transform 1 0 44988 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_482
timestamp 1667941163
transform 1 0 45448 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_490
timestamp 1667941163
transform 1 0 46184 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_514
timestamp 1667941163
transform 1 0 48392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1667941163
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1667941163
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1667941163
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1667941163
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1667941163
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1667941163
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1667941163
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1667941163
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1667941163
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1667941163
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1667941163
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1667941163
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1667941163
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1667941163
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1667941163
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1667941163
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1667941163
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1667941163
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1667941163
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1667941163
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1667941163
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1667941163
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1667941163
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1667941163
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1667941163
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_237
timestamp 1667941163
transform 1 0 22908 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_241
timestamp 1667941163
transform 1 0 23276 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_245
timestamp 1667941163
transform 1 0 23644 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_267
timestamp 1667941163
transform 1 0 25668 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1667941163
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1667941163
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_299
timestamp 1667941163
transform 1 0 28612 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_306
timestamp 1667941163
transform 1 0 29256 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_310
timestamp 1667941163
transform 1 0 29624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_316
timestamp 1667941163
transform 1 0 30176 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_324
timestamp 1667941163
transform 1 0 30912 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_330
timestamp 1667941163
transform 1 0 31464 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1667941163
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_342
timestamp 1667941163
transform 1 0 32568 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_349
timestamp 1667941163
transform 1 0 33212 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_355
timestamp 1667941163
transform 1 0 33764 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_372
timestamp 1667941163
transform 1 0 35328 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_381
timestamp 1667941163
transform 1 0 36156 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_390
timestamp 1667941163
transform 1 0 36984 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_393
timestamp 1667941163
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_400
timestamp 1667941163
transform 1 0 37904 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_407
timestamp 1667941163
transform 1 0 38548 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_419
timestamp 1667941163
transform 1 0 39652 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_426
timestamp 1667941163
transform 1 0 40296 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_438
timestamp 1667941163
transform 1 0 41400 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_446
timestamp 1667941163
transform 1 0 42136 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_449
timestamp 1667941163
transform 1 0 42412 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_467
timestamp 1667941163
transform 1 0 44068 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_479
timestamp 1667941163
transform 1 0 45172 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_491
timestamp 1667941163
transform 1 0 46276 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_502
timestamp 1667941163
transform 1 0 47288 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_505
timestamp 1667941163
transform 1 0 47564 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_510
timestamp 1667941163
transform 1 0 48024 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1667941163
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_8
timestamp 1667941163
transform 1 0 1840 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_15
timestamp 1667941163
transform 1 0 2484 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_22
timestamp 1667941163
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_29
timestamp 1667941163
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_33
timestamp 1667941163
transform 1 0 4140 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_46
timestamp 1667941163
transform 1 0 5336 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_58
timestamp 1667941163
transform 1 0 6440 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_70
timestamp 1667941163
transform 1 0 7544 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1667941163
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1667941163
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1667941163
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1667941163
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1667941163
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1667941163
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1667941163
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1667941163
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1667941163
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1667941163
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1667941163
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1667941163
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1667941163
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1667941163
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1667941163
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1667941163
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_233
timestamp 1667941163
transform 1 0 22540 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_241
timestamp 1667941163
transform 1 0 23276 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_246
timestamp 1667941163
transform 1 0 23736 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1667941163
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1667941163
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_277
timestamp 1667941163
transform 1 0 26588 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_288
timestamp 1667941163
transform 1 0 27600 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_296
timestamp 1667941163
transform 1 0 28336 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_302
timestamp 1667941163
transform 1 0 28888 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1667941163
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_327
timestamp 1667941163
transform 1 0 31188 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_347
timestamp 1667941163
transform 1 0 33028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1667941163
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1667941163
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1667941163
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_370
timestamp 1667941163
transform 1 0 35144 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_376
timestamp 1667941163
transform 1 0 35696 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_393
timestamp 1667941163
transform 1 0 37260 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_405
timestamp 1667941163
transform 1 0 38364 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_417
timestamp 1667941163
transform 1 0 39468 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1667941163
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1667941163
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1667941163
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1667941163
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1667941163
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1667941163
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_477
timestamp 1667941163
transform 1 0 44988 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_485
timestamp 1667941163
transform 1 0 45724 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_489
timestamp 1667941163
transform 1 0 46092 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_514
timestamp 1667941163
transform 1 0 48392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1667941163
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_7
timestamp 1667941163
transform 1 0 1748 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_11
timestamp 1667941163
transform 1 0 2116 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_18
timestamp 1667941163
transform 1 0 2760 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_26
timestamp 1667941163
transform 1 0 3496 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_44
timestamp 1667941163
transform 1 0 5152 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1667941163
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1667941163
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1667941163
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1667941163
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1667941163
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1667941163
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1667941163
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1667941163
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1667941163
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1667941163
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1667941163
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1667941163
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1667941163
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1667941163
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1667941163
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1667941163
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1667941163
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1667941163
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_225
timestamp 1667941163
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_229
timestamp 1667941163
transform 1 0 22172 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_232
timestamp 1667941163
transform 1 0 22448 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_239
timestamp 1667941163
transform 1 0 23092 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_248
timestamp 1667941163
transform 1 0 23920 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_252
timestamp 1667941163
transform 1 0 24288 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_264
timestamp 1667941163
transform 1 0 25392 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1667941163
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_281
timestamp 1667941163
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_286
timestamp 1667941163
transform 1 0 27416 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_294
timestamp 1667941163
transform 1 0 28152 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_313
timestamp 1667941163
transform 1 0 29900 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_320
timestamp 1667941163
transform 1 0 30544 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_332
timestamp 1667941163
transform 1 0 31648 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1667941163
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1667941163
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1667941163
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_373
timestamp 1667941163
transform 1 0 35420 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_379
timestamp 1667941163
transform 1 0 35972 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1667941163
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1667941163
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1667941163
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1667941163
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1667941163
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1667941163
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1667941163
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1667941163
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1667941163
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1667941163
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1667941163
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_497
timestamp 1667941163
transform 1 0 46828 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_502
timestamp 1667941163
transform 1 0 47288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_505
timestamp 1667941163
transform 1 0 47564 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_510
timestamp 1667941163
transform 1 0 48024 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1667941163
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1667941163
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_29
timestamp 1667941163
transform 1 0 3772 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_34
timestamp 1667941163
transform 1 0 4232 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_42
timestamp 1667941163
transform 1 0 4968 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_55
timestamp 1667941163
transform 1 0 6164 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_67
timestamp 1667941163
transform 1 0 7268 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_79
timestamp 1667941163
transform 1 0 8372 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1667941163
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1667941163
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1667941163
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1667941163
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1667941163
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1667941163
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1667941163
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1667941163
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1667941163
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1667941163
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1667941163
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1667941163
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1667941163
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1667941163
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1667941163
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1667941163
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1667941163
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1667941163
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1667941163
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1667941163
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1667941163
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_277
timestamp 1667941163
transform 1 0 26588 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_286
timestamp 1667941163
transform 1 0 27416 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_298
timestamp 1667941163
transform 1 0 28520 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1667941163
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1667941163
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1667941163
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1667941163
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1667941163
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1667941163
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1667941163
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1667941163
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1667941163
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1667941163
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1667941163
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1667941163
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1667941163
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1667941163
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1667941163
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1667941163
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1667941163
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1667941163
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1667941163
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1667941163
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_489
timestamp 1667941163
transform 1 0 46092 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_514
timestamp 1667941163
transform 1 0 48392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1667941163
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_8
timestamp 1667941163
transform 1 0 1840 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_33
timestamp 1667941163
transform 1 0 4140 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1667941163
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1667941163
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_71
timestamp 1667941163
transform 1 0 7636 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_83
timestamp 1667941163
transform 1 0 8740 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_95
timestamp 1667941163
transform 1 0 9844 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_107
timestamp 1667941163
transform 1 0 10948 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1667941163
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1667941163
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1667941163
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1667941163
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1667941163
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1667941163
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1667941163
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1667941163
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1667941163
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1667941163
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1667941163
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1667941163
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1667941163
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1667941163
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1667941163
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1667941163
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1667941163
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1667941163
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1667941163
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1667941163
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1667941163
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1667941163
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1667941163
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1667941163
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1667941163
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1667941163
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1667941163
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1667941163
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1667941163
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1667941163
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1667941163
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1667941163
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1667941163
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1667941163
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1667941163
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1667941163
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1667941163
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1667941163
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1667941163
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1667941163
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_485
timestamp 1667941163
transform 1 0 45724 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_491
timestamp 1667941163
transform 1 0 46276 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_495
timestamp 1667941163
transform 1 0 46644 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_502
timestamp 1667941163
transform 1 0 47288 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_505
timestamp 1667941163
transform 1 0 47564 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_514
timestamp 1667941163
transform 1 0 48392 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1667941163
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_10
timestamp 1667941163
transform 1 0 2024 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1667941163
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_29
timestamp 1667941163
transform 1 0 3772 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_38
timestamp 1667941163
transform 1 0 4600 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_54
timestamp 1667941163
transform 1 0 6072 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_66
timestamp 1667941163
transform 1 0 7176 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_78
timestamp 1667941163
transform 1 0 8280 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1667941163
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1667941163
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1667941163
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1667941163
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1667941163
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1667941163
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1667941163
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1667941163
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1667941163
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1667941163
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1667941163
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1667941163
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1667941163
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1667941163
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1667941163
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1667941163
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1667941163
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1667941163
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1667941163
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1667941163
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1667941163
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1667941163
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1667941163
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1667941163
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1667941163
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1667941163
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1667941163
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1667941163
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1667941163
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1667941163
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1667941163
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1667941163
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1667941163
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1667941163
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1667941163
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1667941163
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_421
timestamp 1667941163
transform 1 0 39836 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_428
timestamp 1667941163
transform 1 0 40480 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_440
timestamp 1667941163
transform 1 0 41584 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_452
timestamp 1667941163
transform 1 0 42688 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_464
timestamp 1667941163
transform 1 0 43792 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_477
timestamp 1667941163
transform 1 0 44988 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_488
timestamp 1667941163
transform 1 0 46000 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_492
timestamp 1667941163
transform 1 0 46368 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_514
timestamp 1667941163
transform 1 0 48392 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1667941163
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_8
timestamp 1667941163
transform 1 0 1840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_33
timestamp 1667941163
transform 1 0 4140 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_49
timestamp 1667941163
transform 1 0 5612 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1667941163
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_57
timestamp 1667941163
transform 1 0 6348 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_62
timestamp 1667941163
transform 1 0 6808 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_74
timestamp 1667941163
transform 1 0 7912 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_86
timestamp 1667941163
transform 1 0 9016 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_98
timestamp 1667941163
transform 1 0 10120 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1667941163
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1667941163
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_113
timestamp 1667941163
transform 1 0 11500 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_121
timestamp 1667941163
transform 1 0 12236 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_125
timestamp 1667941163
transform 1 0 12604 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_132
timestamp 1667941163
transform 1 0 13248 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_157
timestamp 1667941163
transform 1 0 15548 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1667941163
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1667941163
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1667941163
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1667941163
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1667941163
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1667941163
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1667941163
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1667941163
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1667941163
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_249
timestamp 1667941163
transform 1 0 24012 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_256
timestamp 1667941163
transform 1 0 24656 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_265
timestamp 1667941163
transform 1 0 25484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_277
timestamp 1667941163
transform 1 0 26588 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1667941163
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1667941163
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_305
timestamp 1667941163
transform 1 0 29164 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_314
timestamp 1667941163
transform 1 0 29992 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_326
timestamp 1667941163
transform 1 0 31096 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1667941163
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1667941163
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1667941163
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1667941163
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_373
timestamp 1667941163
transform 1 0 35420 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_378
timestamp 1667941163
transform 1 0 35880 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_384
timestamp 1667941163
transform 1 0 36432 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1667941163
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1667941163
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1667941163
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_417
timestamp 1667941163
transform 1 0 39468 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_428
timestamp 1667941163
transform 1 0 40480 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_436
timestamp 1667941163
transform 1 0 41216 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_442
timestamp 1667941163
transform 1 0 41768 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1667941163
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1667941163
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_473
timestamp 1667941163
transform 1 0 44620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_477
timestamp 1667941163
transform 1 0 44988 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_502
timestamp 1667941163
transform 1 0 47288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_505
timestamp 1667941163
transform 1 0 47564 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_510
timestamp 1667941163
transform 1 0 48024 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1667941163
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_26
timestamp 1667941163
transform 1 0 3496 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 1667941163
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_45
timestamp 1667941163
transform 1 0 5244 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_70
timestamp 1667941163
transform 1 0 7544 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1667941163
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1667941163
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1667941163
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_122
timestamp 1667941163
transform 1 0 12328 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_131
timestamp 1667941163
transform 1 0 13156 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1667941163
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_141
timestamp 1667941163
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_164
timestamp 1667941163
transform 1 0 16192 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_171
timestamp 1667941163
transform 1 0 16836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_183
timestamp 1667941163
transform 1 0 17940 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1667941163
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1667941163
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1667941163
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1667941163
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_233
timestamp 1667941163
transform 1 0 22540 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_239
timestamp 1667941163
transform 1 0 23092 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1667941163
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1667941163
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_276
timestamp 1667941163
transform 1 0 26496 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_283
timestamp 1667941163
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_295
timestamp 1667941163
transform 1 0 28244 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1667941163
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1667941163
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_332
timestamp 1667941163
transform 1 0 31648 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_344
timestamp 1667941163
transform 1 0 32752 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_351
timestamp 1667941163
transform 1 0 33396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1667941163
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_365
timestamp 1667941163
transform 1 0 34684 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_373
timestamp 1667941163
transform 1 0 35420 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_395
timestamp 1667941163
transform 1 0 37444 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_399
timestamp 1667941163
transform 1 0 37812 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_403
timestamp 1667941163
transform 1 0 38180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_415
timestamp 1667941163
transform 1 0 39284 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1667941163
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_421
timestamp 1667941163
transform 1 0 39836 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1667941163
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_457
timestamp 1667941163
transform 1 0 43148 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_463
timestamp 1667941163
transform 1 0 43700 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_467
timestamp 1667941163
transform 1 0 44068 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_474
timestamp 1667941163
transform 1 0 44712 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_477
timestamp 1667941163
transform 1 0 44988 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_506
timestamp 1667941163
transform 1 0 47656 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_513
timestamp 1667941163
transform 1 0 48300 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1667941163
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_7
timestamp 1667941163
transform 1 0 1748 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_29
timestamp 1667941163
transform 1 0 3772 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1667941163
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_57
timestamp 1667941163
transform 1 0 6348 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_80
timestamp 1667941163
transform 1 0 8464 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_92
timestamp 1667941163
transform 1 0 9568 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_100
timestamp 1667941163
transform 1 0 10304 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1667941163
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1667941163
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_113
timestamp 1667941163
transform 1 0 11500 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_119
timestamp 1667941163
transform 1 0 12052 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_141
timestamp 1667941163
transform 1 0 14076 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1667941163
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1667941163
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1667941163
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1667941163
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1667941163
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1667941163
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1667941163
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_225
timestamp 1667941163
transform 1 0 21804 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_231
timestamp 1667941163
transform 1 0 22356 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_253
timestamp 1667941163
transform 1 0 24380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1667941163
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1667941163
transform 1 0 26956 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_304
timestamp 1667941163
transform 1 0 29072 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1667941163
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1667941163
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_337
timestamp 1667941163
transform 1 0 32108 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_345
timestamp 1667941163
transform 1 0 32844 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_367
timestamp 1667941163
transform 1 0 34868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_378
timestamp 1667941163
transform 1 0 35880 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_382
timestamp 1667941163
transform 1 0 36248 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_386
timestamp 1667941163
transform 1 0 36616 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1667941163
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_416
timestamp 1667941163
transform 1 0 39376 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1667941163
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1667941163
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1667941163
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_472
timestamp 1667941163
transform 1 0 44528 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_480
timestamp 1667941163
transform 1 0 45264 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_502
timestamp 1667941163
transform 1 0 47288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_505
timestamp 1667941163
transform 1 0 47564 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_510
timestamp 1667941163
transform 1 0 48024 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1667941163
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_12
timestamp 1667941163
transform 1 0 2208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_25
timestamp 1667941163
transform 1 0 3404 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_29
timestamp 1667941163
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_38
timestamp 1667941163
transform 1 0 4600 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_45
timestamp 1667941163
transform 1 0 5244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_52
timestamp 1667941163
transform 1 0 5888 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1667941163
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_62
timestamp 1667941163
transform 1 0 6808 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_69
timestamp 1667941163
transform 1 0 7452 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_76
timestamp 1667941163
transform 1 0 8096 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1667941163
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_90
timestamp 1667941163
transform 1 0 9384 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_102
timestamp 1667941163
transform 1 0 10488 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1667941163
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1667941163
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_121
timestamp 1667941163
transform 1 0 12236 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_125
timestamp 1667941163
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1667941163
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_141
timestamp 1667941163
transform 1 0 14076 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_147
timestamp 1667941163
transform 1 0 14628 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_154
timestamp 1667941163
transform 1 0 15272 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_166
timestamp 1667941163
transform 1 0 16376 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_169
timestamp 1667941163
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_181
timestamp 1667941163
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1667941163
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1667941163
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1667941163
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1667941163
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_225
timestamp 1667941163
transform 1 0 21804 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_233
timestamp 1667941163
transform 1 0 22540 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_239
timestamp 1667941163
transform 1 0 23092 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1667941163
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1667941163
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_264
timestamp 1667941163
transform 1 0 25392 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_276
timestamp 1667941163
transform 1 0 26496 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_281
timestamp 1667941163
transform 1 0 26956 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_286
timestamp 1667941163
transform 1 0 27416 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_293
timestamp 1667941163
transform 1 0 28060 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_301
timestamp 1667941163
transform 1 0 28796 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1667941163
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1667941163
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_314
timestamp 1667941163
transform 1 0 29992 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_326
timestamp 1667941163
transform 1 0 31096 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_334
timestamp 1667941163
transform 1 0 31832 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_337
timestamp 1667941163
transform 1 0 32108 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_345
timestamp 1667941163
transform 1 0 32844 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_350
timestamp 1667941163
transform 1 0 33304 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_362
timestamp 1667941163
transform 1 0 34408 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1667941163
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1667941163
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1667941163
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1667941163
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_401
timestamp 1667941163
transform 1 0 37996 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_405
timestamp 1667941163
transform 1 0 38364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1667941163
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1667941163
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_433
timestamp 1667941163
transform 1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_437
timestamp 1667941163
transform 1 0 41308 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1667941163
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1667941163
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_449
timestamp 1667941163
transform 1 0 42412 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_461
timestamp 1667941163
transform 1 0 43516 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_469
timestamp 1667941163
transform 1 0 44252 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_474
timestamp 1667941163
transform 1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_477
timestamp 1667941163
transform 1 0 44988 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_502
timestamp 1667941163
transform 1 0 47288 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1667941163
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_510
timestamp 1667941163
transform 1 0 48024 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1667941163
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1667941163
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1667941163
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1667941163
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1667941163
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1667941163
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1667941163
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1667941163
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1667941163
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1667941163
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1667941163
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1667941163
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1667941163
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1667941163
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1667941163
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1667941163
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1667941163
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1667941163
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1667941163
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1667941163
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1667941163
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1667941163
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1667941163
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1667941163
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1667941163
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1667941163
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1667941163
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1667941163
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1667941163
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1667941163
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1667941163
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1667941163
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1667941163
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1667941163
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1667941163
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1667941163
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1667941163
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1667941163
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1667941163
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1667941163
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1667941163
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1667941163
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1667941163
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1667941163
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1667941163
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1667941163
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1667941163
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1667941163
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1667941163
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1667941163
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1667941163
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1667941163
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1667941163
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1667941163
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1667941163
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1667941163
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1667941163
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1667941163
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1667941163
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1667941163
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1667941163
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1667941163
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1667941163
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1667941163
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1667941163
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1667941163
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1667941163
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1667941163
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1667941163
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1667941163
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1667941163
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1667941163
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1667941163
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1667941163
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1667941163
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1667941163
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1667941163
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1667941163
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1667941163
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1667941163
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1667941163
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1667941163
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1667941163
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1667941163
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1667941163
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1667941163
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1667941163
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1667941163
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1667941163
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1667941163
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1667941163
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1667941163
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1667941163
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1667941163
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1667941163
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1667941163
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1667941163
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1667941163
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1667941163
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1667941163
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1667941163
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1667941163
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1667941163
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1667941163
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1667941163
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1667941163
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1667941163
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1667941163
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1667941163
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1667941163
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1667941163
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1667941163
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1667941163
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1667941163
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1667941163
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1667941163
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1667941163
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1667941163
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1667941163
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1667941163
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1667941163
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1667941163
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1667941163
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1667941163
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1667941163
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1667941163
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1667941163
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1667941163
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1667941163
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1667941163
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1667941163
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1667941163
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1667941163
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1667941163
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1667941163
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1667941163
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1667941163
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1667941163
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1667941163
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1667941163
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1667941163
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1667941163
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1667941163
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1667941163
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1667941163
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1667941163
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1667941163
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1667941163
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1667941163
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1667941163
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1667941163
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1667941163
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1667941163
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1667941163
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1667941163
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1667941163
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1667941163
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1667941163
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1667941163
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1667941163
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1667941163
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1667941163
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1667941163
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1667941163
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1667941163
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1667941163
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1667941163
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1667941163
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1667941163
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1667941163
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1667941163
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1667941163
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1667941163
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1667941163
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1667941163
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1667941163
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1667941163
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1667941163
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1667941163
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1667941163
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1667941163
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1667941163
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1667941163
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1667941163
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1667941163
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1667941163
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1667941163
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1667941163
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1667941163
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1667941163
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1667941163
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1667941163
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1667941163
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1667941163
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1667941163
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1667941163
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1667941163
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1667941163
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1667941163
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1667941163
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1667941163
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1667941163
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1667941163
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1667941163
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1667941163
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1667941163
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1667941163
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1667941163
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1667941163
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1667941163
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1667941163
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1667941163
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1667941163
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1667941163
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1667941163
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1667941163
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1667941163
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1667941163
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1667941163
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1667941163
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1667941163
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1667941163
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1667941163
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1667941163
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1667941163
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1667941163
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1667941163
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1667941163
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1667941163
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1667941163
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1667941163
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1667941163
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1667941163
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1667941163
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1667941163
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1667941163
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1667941163
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1667941163
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1667941163
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1667941163
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1667941163
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1667941163
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1667941163
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _0663_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2576 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _0664_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  _0665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 1748 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 45724 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 47748 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 47012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 47012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 47748 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0676_
timestamp 1667941163
transform 1 0 41032 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 4324 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 45172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 26864 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 47748 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 47748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 6532 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 47012 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0687_
timestamp 1667941163
transform 1 0 4140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 47748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 29716 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 47012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 47012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 1932 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 2484 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 47748 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0698_
timestamp 1667941163
transform 1 0 2392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 33120 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 22816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 44436 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 48024 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 47012 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 5520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 47748 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0709_
timestamp 1667941163
transform 1 0 4508 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 40664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 46736 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 28336 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 45632 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 45816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 45816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 40204 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0720_
timestamp 1667941163
transform 1 0 4232 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 2300 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 32292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 37904 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 36524 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0731_
timestamp 1667941163
transform 1 0 4968 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 5612 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 47748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 47748 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 47748 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 16560 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 46368 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 39284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 41492 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 12328 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0742_
timestamp 1667941163
transform 1 0 6532 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 47748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 2760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 2300 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 47748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 46368 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 47748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 47012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 12972 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0753_
timestamp 1667941163
transform 1 0 5060 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 43700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 35604 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 13524 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 47748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 25208 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 47748 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 24380 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 28980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0764_
timestamp 1667941163
transform 1 0 4508 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 42780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 1564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 47748 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 3956 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 41308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 2300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 44436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 10488 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 2760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 44344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 47012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 47012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 2576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 47012 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 43332 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 45080 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 41860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 38916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 36432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 36708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0789_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36156 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 36984 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0792_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37260 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 37628 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0794_
timestamp 1667941163
transform 1 0 36248 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0795_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35972 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0797_
timestamp 1667941163
transform 1 0 37536 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0798_
timestamp 1667941163
transform 1 0 37352 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0799_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38916 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0800_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 41400 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0801_
timestamp 1667941163
transform 1 0 43792 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 45908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0803_
timestamp 1667941163
transform 1 0 33580 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 44160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 26404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 26128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 25208 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 27416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0811_
timestamp 1667941163
transform 1 0 27232 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 28060 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 28612 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0814_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28428 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0815_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0816_
timestamp 1667941163
transform 1 0 27600 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0817_
timestamp 1667941163
transform 1 0 27416 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0818_
timestamp 1667941163
transform 1 0 26312 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0819_
timestamp 1667941163
transform 1 0 27140 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0820_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0821_
timestamp 1667941163
transform 1 0 27140 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0822_
timestamp 1667941163
transform 1 0 27324 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0823_
timestamp 1667941163
transform 1 0 32292 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_1  _0824_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26956 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 30360 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0826_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0827_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 46000 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 46276 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 45632 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 43976 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 43792 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 41860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0834_
timestamp 1667941163
transform 1 0 42504 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 40664 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 40020 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0837_
timestamp 1667941163
transform 1 0 40020 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 37444 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38916 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38824 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0841_
timestamp 1667941163
transform 1 0 39560 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0842_
timestamp 1667941163
transform 1 0 40572 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0843_
timestamp 1667941163
transform 1 0 40296 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1667941163
transform 1 0 43516 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0845_
timestamp 1667941163
transform 1 0 42872 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0846_
timestamp 1667941163
transform 1 0 44804 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0847_
timestamp 1667941163
transform 1 0 45172 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 45448 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0849_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 46092 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0850_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33672 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35236 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0853_
timestamp 1667941163
transform 1 0 34868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0854_
timestamp 1667941163
transform 1 0 34868 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0856_
timestamp 1667941163
transform 1 0 37444 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0857_
timestamp 1667941163
transform 1 0 37720 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0858_
timestamp 1667941163
transform 1 0 37444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0859_
timestamp 1667941163
transform 1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0860_
timestamp 1667941163
transform 1 0 38732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0861_
timestamp 1667941163
transform 1 0 38640 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0862_
timestamp 1667941163
transform 1 0 40020 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0863_
timestamp 1667941163
transform 1 0 39928 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0864_
timestamp 1667941163
transform 1 0 40756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1667941163
transform 1 0 41584 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0866_
timestamp 1667941163
transform 1 0 40848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0867_
timestamp 1667941163
transform 1 0 42136 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1667941163
transform 1 0 41400 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0869_
timestamp 1667941163
transform 1 0 42044 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0870_
timestamp 1667941163
transform 1 0 31556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0871_
timestamp 1667941163
transform 1 0 29808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0872_
timestamp 1667941163
transform 1 0 29716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0873_
timestamp 1667941163
transform 1 0 31188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0874_
timestamp 1667941163
transform 1 0 30912 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0875_
timestamp 1667941163
transform 1 0 30544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0876_
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0877_
timestamp 1667941163
transform 1 0 32292 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1667941163
transform 1 0 33028 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0879_
timestamp 1667941163
transform 1 0 30636 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0880_
timestamp 1667941163
transform 1 0 30912 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1667941163
transform 1 0 29992 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0882_
timestamp 1667941163
transform 1 0 30728 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0883_
timestamp 1667941163
transform 1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0884_
timestamp 1667941163
transform 1 0 29808 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 1667941163
transform 1 0 29808 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0886_
timestamp 1667941163
transform 1 0 31556 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0888_
timestamp 1667941163
transform 1 0 30360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0889_
timestamp 1667941163
transform 1 0 29440 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0890_
timestamp 1667941163
transform 1 0 37904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0891_
timestamp 1667941163
transform 1 0 39192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0892_
timestamp 1667941163
transform 1 0 40020 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0893_
timestamp 1667941163
transform 1 0 40020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0894_
timestamp 1667941163
transform 1 0 40020 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0895_
timestamp 1667941163
transform 1 0 39100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0896_
timestamp 1667941163
transform 1 0 41676 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0897_
timestamp 1667941163
transform 1 0 41492 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0898_
timestamp 1667941163
transform 1 0 42228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0899_
timestamp 1667941163
transform 1 0 44344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0900_
timestamp 1667941163
transform 1 0 43424 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0901_
timestamp 1667941163
transform 1 0 43332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0902_
timestamp 1667941163
transform 1 0 43700 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0903_
timestamp 1667941163
transform 1 0 42964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1667941163
transform 1 0 45724 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0905_
timestamp 1667941163
transform 1 0 46552 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1667941163
transform 1 0 46368 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0907_
timestamp 1667941163
transform 1 0 45632 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0908_
timestamp 1667941163
transform 1 0 45540 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1667941163
transform 1 0 33396 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0910_
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36156 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0912_
timestamp 1667941163
transform 1 0 34224 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1667941163
transform 1 0 35972 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1667941163
transform 1 0 35328 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34960 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0916_
timestamp 1667941163
transform 1 0 38180 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0917_
timestamp 1667941163
transform 1 0 34776 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0918_
timestamp 1667941163
transform 1 0 33488 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0919_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0920_
timestamp 1667941163
transform 1 0 36340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0921_
timestamp 1667941163
transform 1 0 35420 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1667941163
transform 1 0 36340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0923_
timestamp 1667941163
transform 1 0 35144 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0924_
timestamp 1667941163
transform 1 0 35512 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0925_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35144 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0926_
timestamp 1667941163
transform 1 0 37444 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 41124 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0929_
timestamp 1667941163
transform 1 0 35144 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1667941163
transform 1 0 34868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0931_
timestamp 1667941163
transform 1 0 34868 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0932_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35880 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0933_
timestamp 1667941163
transform 1 0 32844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0935_
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0936_
timestamp 1667941163
transform 1 0 34132 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0937_
timestamp 1667941163
transform 1 0 35236 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0939_
timestamp 1667941163
transform 1 0 34868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0940_
timestamp 1667941163
transform 1 0 35788 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0941_
timestamp 1667941163
transform 1 0 37720 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0942_
timestamp 1667941163
transform 1 0 34592 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0943_
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34868 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0945_
timestamp 1667941163
transform 1 0 37536 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0946_
timestamp 1667941163
transform 1 0 38548 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0947_
timestamp 1667941163
transform 1 0 38456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0948_
timestamp 1667941163
transform 1 0 37904 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0949_
timestamp 1667941163
transform 1 0 37812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0950_
timestamp 1667941163
transform 1 0 39836 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0951_
timestamp 1667941163
transform 1 0 39008 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0952_
timestamp 1667941163
transform 1 0 40020 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1667941163
transform 1 0 41124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0954_
timestamp 1667941163
transform 1 0 40940 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0955_
timestamp 1667941163
transform 1 0 44068 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1667941163
transform 1 0 43792 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1667941163
transform 1 0 43792 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0958_
timestamp 1667941163
transform 1 0 40020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0959_
timestamp 1667941163
transform 1 0 40112 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0960_
timestamp 1667941163
transform 1 0 43148 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0961_
timestamp 1667941163
transform 1 0 43148 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0962_
timestamp 1667941163
transform 1 0 42964 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0963_
timestamp 1667941163
transform 1 0 44160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0964_
timestamp 1667941163
transform 1 0 43700 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0965_
timestamp 1667941163
transform 1 0 43884 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0966_
timestamp 1667941163
transform 1 0 40940 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0967_
timestamp 1667941163
transform 1 0 41584 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0968_
timestamp 1667941163
transform 1 0 36432 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0969_
timestamp 1667941163
transform 1 0 24840 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1667941163
transform 1 0 24196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0971_
timestamp 1667941163
transform 1 0 34868 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1667941163
transform 1 0 35880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0973_
timestamp 1667941163
transform 1 0 26404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0974_
timestamp 1667941163
transform 1 0 27140 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0975_
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0976_
timestamp 1667941163
transform 1 0 27048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0977_
timestamp 1667941163
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0978_
timestamp 1667941163
transform 1 0 22632 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0979_
timestamp 1667941163
transform 1 0 29716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0980_
timestamp 1667941163
transform 1 0 30544 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0981_
timestamp 1667941163
transform 1 0 25944 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0982_
timestamp 1667941163
transform 1 0 26128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0983_
timestamp 1667941163
transform 1 0 26128 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 1667941163
transform 1 0 26036 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0985_
timestamp 1667941163
transform 1 0 27140 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0986_
timestamp 1667941163
transform 1 0 26404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0987_
timestamp 1667941163
transform 1 0 26680 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0989_
timestamp 1667941163
transform 1 0 27140 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0990_
timestamp 1667941163
transform 1 0 26312 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0991_
timestamp 1667941163
transform 1 0 26128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0992_
timestamp 1667941163
transform 1 0 25852 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0994_
timestamp 1667941163
transform 1 0 24380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0995_
timestamp 1667941163
transform 1 0 23276 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0996_
timestamp 1667941163
transform 1 0 23368 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0997_
timestamp 1667941163
transform 1 0 23276 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0998_
timestamp 1667941163
transform 1 0 26404 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0999_
timestamp 1667941163
transform 1 0 24840 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1000_
timestamp 1667941163
transform 1 0 23000 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 1667941163
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1002_
timestamp 1667941163
transform 1 0 23644 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1003_
timestamp 1667941163
transform 1 0 22724 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1004_
timestamp 1667941163
transform 1 0 23276 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1005_
timestamp 1667941163
transform 1 0 22080 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1667941163
transform 1 0 22356 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1008_
timestamp 1667941163
transform 1 0 23000 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1667941163
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1010_
timestamp 1667941163
transform 1 0 22080 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1011_
timestamp 1667941163
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1012_
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1014_
timestamp 1667941163
transform 1 0 25208 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1015_
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1016_
timestamp 1667941163
transform 1 0 22448 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1017_
timestamp 1667941163
transform 1 0 23184 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1018_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1019_
timestamp 1667941163
transform 1 0 23092 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1020_
timestamp 1667941163
transform 1 0 22908 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1021_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1667941163
transform 1 0 23276 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1023_
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1024_
timestamp 1667941163
transform 1 0 25852 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1025_
timestamp 1667941163
transform 1 0 26036 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1026_
timestamp 1667941163
transform 1 0 27508 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1027_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1028_
timestamp 1667941163
transform 1 0 36892 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 36708 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1667941163
transform 1 0 27140 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 27140 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1032_
timestamp 1667941163
transform 1 0 40020 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1033_
timestamp 1667941163
transform 1 0 38824 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1034_
timestamp 1667941163
transform 1 0 41216 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1035_
timestamp 1667941163
transform 1 0 40940 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1036_
timestamp 1667941163
transform 1 0 38272 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38548 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1038_
timestamp 1667941163
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1039_
timestamp 1667941163
transform 1 0 38272 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1040_
timestamp 1667941163
transform 1 0 37444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1041_
timestamp 1667941163
transform 1 0 40020 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1042_
timestamp 1667941163
transform 1 0 40020 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1043_
timestamp 1667941163
transform 1 0 40756 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1044_
timestamp 1667941163
transform 1 0 40664 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1045_
timestamp 1667941163
transform 1 0 39284 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1667941163
transform 1 0 40020 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1047_
timestamp 1667941163
transform 1 0 38180 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1048_
timestamp 1667941163
transform 1 0 38548 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1049_
timestamp 1667941163
transform 1 0 38548 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1050_
timestamp 1667941163
transform 1 0 37444 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1051_
timestamp 1667941163
transform 1 0 40480 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1052_
timestamp 1667941163
transform 1 0 39284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38732 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1667941163
transform 1 0 40020 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1055_
timestamp 1667941163
transform 1 0 39284 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1056_
timestamp 1667941163
transform 1 0 38916 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1057_
timestamp 1667941163
transform 1 0 38088 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1058_
timestamp 1667941163
transform 1 0 42596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1059_
timestamp 1667941163
transform 1 0 40388 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1060_
timestamp 1667941163
transform 1 0 40756 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1061_
timestamp 1667941163
transform 1 0 40848 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1062_
timestamp 1667941163
transform 1 0 40940 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1063_
timestamp 1667941163
transform 1 0 40756 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1064_
timestamp 1667941163
transform 1 0 39928 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1065_
timestamp 1667941163
transform 1 0 43332 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1667941163
transform 1 0 43884 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1067_
timestamp 1667941163
transform 1 0 44344 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1068_
timestamp 1667941163
transform 1 0 43424 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1069_
timestamp 1667941163
transform 1 0 42872 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1070_
timestamp 1667941163
transform 1 0 45080 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1071_
timestamp 1667941163
transform 1 0 44804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1072_
timestamp 1667941163
transform 1 0 45908 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1073_
timestamp 1667941163
transform 1 0 46920 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1074_
timestamp 1667941163
transform 1 0 46828 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1075_
timestamp 1667941163
transform 1 0 43976 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1076_
timestamp 1667941163
transform 1 0 44620 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1077_
timestamp 1667941163
transform 1 0 44068 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1078_
timestamp 1667941163
transform 1 0 45172 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1079_
timestamp 1667941163
transform 1 0 45172 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1080_
timestamp 1667941163
transform 1 0 43976 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1667941163
transform 1 0 43148 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1667941163
transform 1 0 42872 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1083_
timestamp 1667941163
transform 1 0 44068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1084_
timestamp 1667941163
transform 1 0 45356 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1085_
timestamp 1667941163
transform 1 0 45632 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1086_
timestamp 1667941163
transform 1 0 46828 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1087_
timestamp 1667941163
transform 1 0 46644 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1088_
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1667941163
transform 1 0 24840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1090_
timestamp 1667941163
transform 1 0 33396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1091_
timestamp 1667941163
transform 1 0 29716 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1667941163
transform 1 0 28704 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1093_
timestamp 1667941163
transform 1 0 31188 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1667941163
transform 1 0 31464 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1095_
timestamp 1667941163
transform 1 0 32292 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1096_
timestamp 1667941163
transform 1 0 33120 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1097_
timestamp 1667941163
transform 1 0 30176 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1667941163
transform 1 0 29716 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1099_
timestamp 1667941163
transform 1 0 29716 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1100_
timestamp 1667941163
transform 1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1101_
timestamp 1667941163
transform 1 0 29716 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1667941163
transform 1 0 28980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 1667941163
transform 1 0 30544 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1104_
timestamp 1667941163
transform 1 0 31372 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1105_
timestamp 1667941163
transform 1 0 38824 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1667941163
transform 1 0 40020 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30912 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1108_
timestamp 1667941163
transform 1 0 32292 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31280 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1110_
timestamp 1667941163
transform 1 0 30912 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1667941163
transform 1 0 31280 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1113_
timestamp 1667941163
transform 1 0 39836 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1667941163
transform 1 0 40020 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1115_
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1667941163
transform 1 0 35880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1117_
timestamp 1667941163
transform 1 0 33672 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1118_
timestamp 1667941163
transform 1 0 34132 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1119_
timestamp 1667941163
transform 1 0 34868 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1120_
timestamp 1667941163
transform 1 0 35696 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1121_
timestamp 1667941163
transform 1 0 33120 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1667941163
transform 1 0 32476 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1667941163
transform 1 0 33028 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1124_
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1125_
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1126_
timestamp 1667941163
transform 1 0 31004 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1127_
timestamp 1667941163
transform 1 0 31004 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1128_
timestamp 1667941163
transform 1 0 32660 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1667941163
transform 1 0 33488 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1130_
timestamp 1667941163
transform 1 0 33028 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 1667941163
transform 1 0 34500 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1133_
timestamp 1667941163
transform 1 0 33120 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36156 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1135_
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1136_
timestamp 1667941163
transform 1 0 22632 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1137_
timestamp 1667941163
transform 1 0 23460 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 1667941163
transform 1 0 27968 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1139_
timestamp 1667941163
transform 1 0 28244 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1140_
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1667941163
transform 1 0 23184 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1142_
timestamp 1667941163
transform 1 0 24104 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1143_
timestamp 1667941163
transform 1 0 23828 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1145_
timestamp 1667941163
transform 1 0 24564 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1146_
timestamp 1667941163
transform 1 0 24564 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1667941163
transform 1 0 23828 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1148_
timestamp 1667941163
transform 1 0 24564 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1667941163
transform 1 0 23828 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1150_
timestamp 1667941163
transform 1 0 25576 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1151_
timestamp 1667941163
transform 1 0 26404 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1152_
timestamp 1667941163
transform 1 0 25392 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1153_
timestamp 1667941163
transform 1 0 24932 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1154_
timestamp 1667941163
transform 1 0 27140 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1155_
timestamp 1667941163
transform 1 0 25484 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1156_
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1157_
timestamp 1667941163
transform 1 0 25760 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 1667941163
transform 1 0 26956 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1159_
timestamp 1667941163
transform 1 0 27140 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1160_
timestamp 1667941163
transform 1 0 27416 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1161_
timestamp 1667941163
transform 1 0 28520 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1667941163
transform 1 0 29716 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1163_
timestamp 1667941163
transform 1 0 27968 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1164_
timestamp 1667941163
transform 1 0 36616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1165_
timestamp 1667941163
transform 1 0 28520 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1166_
timestamp 1667941163
transform 1 0 27324 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1167_
timestamp 1667941163
transform 1 0 28428 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1168_
timestamp 1667941163
transform 1 0 28980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1169_
timestamp 1667941163
transform 1 0 29716 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1170_
timestamp 1667941163
transform 1 0 30268 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 1667941163
transform 1 0 31004 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1667941163
transform 1 0 32936 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1173_
timestamp 1667941163
transform 1 0 32292 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1667941163
transform 1 0 32292 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1175_
timestamp 1667941163
transform 1 0 30544 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1176_
timestamp 1667941163
transform 1 0 29716 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1177_
timestamp 1667941163
transform 1 0 28520 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1178_
timestamp 1667941163
transform 1 0 30544 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1179_
timestamp 1667941163
transform 1 0 30452 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1180_
timestamp 1667941163
transform 1 0 28244 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1181_
timestamp 1667941163
transform -1 0 23920 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1182_
timestamp 1667941163
transform 1 0 23368 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1183_
timestamp 1667941163
transform 1 0 31924 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1184_
timestamp 1667941163
transform 1 0 32844 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1185_
timestamp 1667941163
transform 1 0 33856 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1667941163
transform 1 0 33764 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1667941163
transform 1 0 34868 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1667941163
transform 1 0 34868 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1667941163
transform 1 0 35696 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1667941163
transform 1 0 35696 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1191_
timestamp 1667941163
transform 1 0 37444 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1192_
timestamp 1667941163
transform 1 0 36708 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1193_
timestamp 1667941163
transform 1 0 38180 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1194_
timestamp 1667941163
transform 1 0 38272 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1195_
timestamp 1667941163
transform 1 0 40020 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1196_
timestamp 1667941163
transform 1 0 39192 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1197_
timestamp 1667941163
transform 1 0 36892 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1198_
timestamp 1667941163
transform 1 0 35512 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1199_
timestamp 1667941163
transform 1 0 35052 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1200_
timestamp 1667941163
transform 1 0 36432 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1201_
timestamp 1667941163
transform 1 0 36248 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1202_
timestamp 1667941163
transform 1 0 35144 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1667941163
transform 1 0 41492 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1204_
timestamp 1667941163
transform 1 0 42596 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 1667941163
transform 1 0 43884 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1667941163
transform 1 0 43056 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1207_
timestamp 1667941163
transform 1 0 45172 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1667941163
transform 1 0 45172 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1209_
timestamp 1667941163
transform 1 0 43884 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1667941163
transform 1 0 45172 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1211_
timestamp 1667941163
transform 1 0 45172 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1667941163
transform 1 0 45172 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1213_
timestamp 1667941163
transform 1 0 42688 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1667941163
transform 1 0 43516 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1215_
timestamp 1667941163
transform 1 0 41400 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1216_
timestamp 1667941163
transform 1 0 41032 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1217_
timestamp 1667941163
transform 1 0 41676 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1218_
timestamp 1667941163
transform 1 0 42320 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1219_
timestamp 1667941163
transform 1 0 42596 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1220_
timestamp 1667941163
transform 1 0 44068 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1221_
timestamp 1667941163
transform 1 0 44160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1222_
timestamp 1667941163
transform 1 0 42780 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1667941163
transform 1 0 43332 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1224_
timestamp 1667941163
transform 1 0 42504 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32936 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1226_
timestamp 1667941163
transform 1 0 33396 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1227_
timestamp 1667941163
transform 1 0 33580 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1228_
timestamp 1667941163
transform 1 0 37260 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1229_
timestamp 1667941163
transform 1 0 38456 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1230_
timestamp 1667941163
transform 1 0 40112 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1231_
timestamp 1667941163
transform 1 0 42596 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1232_
timestamp 1667941163
transform 1 0 43240 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 1667941163
transform 1 0 31556 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1667941163
transform 1 0 31280 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 1667941163
transform 1 0 31188 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1667941163
transform 1 0 29900 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 1667941163
transform 1 0 29716 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1667941163
transform 1 0 29716 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1667941163
transform 1 0 37444 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1667941163
transform 1 0 39100 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1667941163
transform 1 0 38548 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1667941163
transform 1 0 40664 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1667941163
transform 1 0 43240 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1667941163
transform 1 0 42872 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1667941163
transform 1 0 45816 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1667941163
transform 1 0 45540 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1667941163
transform 1 0 34040 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1667941163
transform 1 0 32936 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1667941163
transform 1 0 35512 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1667941163
transform 1 0 32292 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1667941163
transform 1 0 34868 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1667941163
transform 1 0 37720 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1667941163
transform 1 0 40480 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1667941163
transform 1 0 43240 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1667941163
transform 1 0 41584 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1667941163
transform 1 0 34868 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1667941163
transform 1 0 28704 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1667941163
transform 1 0 27232 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1667941163
transform 1 0 24656 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1667941163
transform 1 0 24380 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1667941163
transform 1 0 26864 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1667941163
transform 1 0 37444 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1667941163
transform 1 0 26036 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1667941163
transform 1 0 36340 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1667941163
transform 1 0 36708 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1667941163
transform 1 0 37444 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1667941163
transform 1 0 41492 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1667941163
transform 1 0 42964 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1667941163
transform 1 0 46920 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1667941163
transform 1 0 42780 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1667941163
transform 1 0 46920 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1667941163
transform 1 0 27784 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1667941163
transform 1 0 29348 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp 1667941163
transform 1 0 31280 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1667941163
transform 1 0 32200 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1667941163
transform 1 0 28704 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1667941163
transform 1 0 28244 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1667941163
transform 1 0 30360 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1667941163
transform 1 0 39652 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1667941163
transform 1 0 32108 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1667941163
transform 1 0 38088 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1667941163
transform 1 0 35420 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1667941163
transform 1 0 34224 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1667941163
transform 1 0 34500 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1667941163
transform 1 0 32292 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1667941163
transform 1 0 30268 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1667941163
transform 1 0 30820 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1667941163
transform 1 0 32568 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1667941163
transform 1 0 24196 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1667941163
transform 1 0 27140 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1667941163
transform 1 0 24564 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1667941163
transform 1 0 23920 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1667941163
transform 1 0 23552 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1667941163
transform 1 0 23644 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1667941163
transform 1 0 24196 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1667941163
transform 1 0 25484 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1667941163
transform 1 0 25576 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1667941163
transform 1 0 27140 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1667941163
transform 1 0 28060 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1667941163
transform 1 0 28612 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1667941163
transform 1 0 26680 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1667941163
transform 1 0 28428 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1311_
timestamp 1667941163
transform 1 0 29716 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp 1667941163
transform 1 0 31556 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp 1667941163
transform 1 0 31556 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp 1667941163
transform 1 0 28060 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1667941163
transform 1 0 24564 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1667941163
transform 1 0 33120 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1667941163
transform 1 0 32936 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1667941163
transform 1 0 33856 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1667941163
transform 1 0 35788 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1667941163
transform 1 0 36340 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1667941163
transform 1 0 38180 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1667941163
transform 1 0 38640 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1667941163
transform 1 0 35420 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1667941163
transform 1 0 42044 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1667941163
transform 1 0 43700 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1667941163
transform 1 0 45816 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1667941163
transform 1 0 44712 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1667941163
transform 1 0 44620 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1667941163
transform 1 0 42596 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1667941163
transform 1 0 40848 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1667941163
transform 1 0 42688 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1667941163
transform 1 0 40664 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1437__9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7544 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1438__10
timestamp 1667941163
transform 1 0 1564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1438_
timestamp 1667941163
transform 1 0 2208 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1439__11
timestamp 1667941163
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1439_
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1440__12
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1440_
timestamp 1667941163
transform 1 0 2116 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1441__13
timestamp 1667941163
transform 1 0 43700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1441_
timestamp 1667941163
transform 1 0 45172 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1442_
timestamp 1667941163
transform 1 0 3772 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1442__14
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1443__15
timestamp 1667941163
transform 1 0 47748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1443_
timestamp 1667941163
transform 1 0 46460 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1444__16
timestamp 1667941163
transform 1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1444_
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1445__17
timestamp 1667941163
transform 1 0 47748 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1445_
timestamp 1667941163
transform 1 0 46460 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1446__18
timestamp 1667941163
transform 1 0 47748 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1446_
timestamp 1667941163
transform 1 0 45724 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1447__19
timestamp 1667941163
transform 1 0 47748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1447_
timestamp 1667941163
transform 1 0 46460 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1448__20
timestamp 1667941163
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1448_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1449_
timestamp 1667941163
transform 1 0 45356 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1449__21
timestamp 1667941163
transform 1 0 44712 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1450__22
timestamp 1667941163
transform 1 0 4324 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1450_
timestamp 1667941163
transform 1 0 4140 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1451__23
timestamp 1667941163
transform 1 0 27140 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1451_
timestamp 1667941163
transform 1 0 27140 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1452__24
timestamp 1667941163
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1452_
timestamp 1667941163
transform 1 0 1840 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1453__25
timestamp 1667941163
transform 1 0 47012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1453_
timestamp 1667941163
transform 1 0 46460 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1454__26
timestamp 1667941163
transform 1 0 47012 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1454_
timestamp 1667941163
transform 1 0 46460 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1455__27
timestamp 1667941163
transform 1 0 4968 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1455_
timestamp 1667941163
transform 1 0 5612 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1456_
timestamp 1667941163
transform 1 0 45356 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1456__28
timestamp 1667941163
transform 1 0 47748 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1457__29
timestamp 1667941163
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1457_
timestamp 1667941163
transform 1 0 2116 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1458__30
timestamp 1667941163
transform 1 0 45816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1458_
timestamp 1667941163
transform 1 0 46460 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1459__31
timestamp 1667941163
transform 1 0 29716 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1459_
timestamp 1667941163
transform 1 0 29716 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1460__32
timestamp 1667941163
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1460_
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1461__33
timestamp 1667941163
transform 1 0 47748 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1461_
timestamp 1667941163
transform 1 0 46460 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1462_
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1462__34
timestamp 1667941163
transform 1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1463_
timestamp 1667941163
transform 1 0 46460 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1463__35
timestamp 1667941163
transform 1 0 47748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1464_
timestamp 1667941163
transform 1 0 1564 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1464__36
timestamp 1667941163
transform 1 0 2852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1465__37
timestamp 1667941163
transform 1 0 44344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1465_
timestamp 1667941163
transform 1 0 44896 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1466_
timestamp 1667941163
transform 1 0 6164 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1466__38
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1467__39
timestamp 1667941163
transform 1 0 47748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1467_
timestamp 1667941163
transform 1 0 46460 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1468_
timestamp 1667941163
transform 1 0 45356 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1468__40
timestamp 1667941163
transform 1 0 43792 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1469__41
timestamp 1667941163
transform 1 0 47012 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1469_
timestamp 1667941163
transform 1 0 46460 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1470__42
timestamp 1667941163
transform 1 0 33028 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1470_
timestamp 1667941163
transform 1 0 32936 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1471_
timestamp 1667941163
transform 1 0 6716 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1471__43
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1472_
timestamp 1667941163
transform 1 0 1564 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1472__44
timestamp 1667941163
transform 1 0 1840 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1473__45
timestamp 1667941163
transform 1 0 47012 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1473_
timestamp 1667941163
transform 1 0 46460 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1474__46
timestamp 1667941163
transform 1 0 22816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1474_
timestamp 1667941163
transform 1 0 22448 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1475__47
timestamp 1667941163
transform 1 0 44436 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1475_
timestamp 1667941163
transform 1 0 45356 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1476__48
timestamp 1667941163
transform 1 0 2116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1476_
timestamp 1667941163
transform 1 0 2024 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1477__49
timestamp 1667941163
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1477_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1478__50
timestamp 1667941163
transform 1 0 1748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1478_
timestamp 1667941163
transform 1 0 2024 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1479_
timestamp 1667941163
transform 1 0 46460 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1479__51
timestamp 1667941163
transform 1 0 47748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1480__52
timestamp 1667941163
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1480_
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1481_
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1481__53
timestamp 1667941163
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1482__54
timestamp 1667941163
transform 1 0 40020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1482_
timestamp 1667941163
transform 1 0 40020 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1483_
timestamp 1667941163
transform 1 0 46460 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1484_
timestamp 1667941163
transform 1 0 27692 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1485_
timestamp 1667941163
transform 1 0 45356 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1486_
timestamp 1667941163
transform 1 0 45908 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1487__55
timestamp 1667941163
transform 1 0 47932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1487_
timestamp 1667941163
transform 1 0 45632 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1488__56
timestamp 1667941163
transform 1 0 2116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1488_
timestamp 1667941163
transform 1 0 2024 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1489__57
timestamp 1667941163
transform 1 0 40204 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1489_
timestamp 1667941163
transform 1 0 40112 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1490__58
timestamp 1667941163
transform 1 0 2116 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1490_
timestamp 1667941163
transform 1 0 2024 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1491__59
timestamp 1667941163
transform 1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1491_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1492_
timestamp 1667941163
transform 1 0 46460 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1492__60
timestamp 1667941163
transform 1 0 47748 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1493__61
timestamp 1667941163
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1493_
timestamp 1667941163
transform 1 0 27416 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1494_
timestamp 1667941163
transform 1 0 37444 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1494__62
timestamp 1667941163
transform 1 0 36340 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1495__63
timestamp 1667941163
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1495_
timestamp 1667941163
transform 1 0 2116 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1496__64
timestamp 1667941163
transform 1 0 38088 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1496_
timestamp 1667941163
transform 1 0 39744 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1497__65
timestamp 1667941163
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1497_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1498__66
timestamp 1667941163
transform 1 0 38640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1498_
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1499_
timestamp 1667941163
transform 1 0 2024 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1499__67
timestamp 1667941163
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1500_
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1500__68
timestamp 1667941163
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1501__69
timestamp 1667941163
transform 1 0 6532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1501_
timestamp 1667941163
transform 1 0 6532 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1502__70
timestamp 1667941163
transform 1 0 47748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1502_
timestamp 1667941163
transform 1 0 46460 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1503__71
timestamp 1667941163
transform 1 0 47012 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1503_
timestamp 1667941163
transform 1 0 46460 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1504__72
timestamp 1667941163
transform 1 0 47012 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1504_
timestamp 1667941163
transform 1 0 46460 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1505__73
timestamp 1667941163
transform 1 0 14996 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1505_
timestamp 1667941163
transform 1 0 14444 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1506__74
timestamp 1667941163
transform 1 0 47748 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1506_
timestamp 1667941163
transform 1 0 46460 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1507__75
timestamp 1667941163
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1507_
timestamp 1667941163
transform 1 0 25852 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1508_
timestamp 1667941163
transform 1 0 38640 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1508__76
timestamp 1667941163
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1509__77
timestamp 1667941163
transform 1 0 41400 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1509_
timestamp 1667941163
transform 1 0 42596 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1510__78
timestamp 1667941163
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1510_
timestamp 1667941163
transform 1 0 24748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1511_
timestamp 1667941163
transform 1 0 46460 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1511__79
timestamp 1667941163
transform 1 0 47748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1512__80
timestamp 1667941163
transform 1 0 2116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1512_
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1513_
timestamp 1667941163
transform 1 0 46460 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1513__81
timestamp 1667941163
transform 1 0 47748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1514__82
timestamp 1667941163
transform 1 0 12328 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1514_
timestamp 1667941163
transform 1 0 12144 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1515__83
timestamp 1667941163
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1515_
timestamp 1667941163
transform 1 0 4692 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1516_
timestamp 1667941163
transform 1 0 10304 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1516__84
timestamp 1667941163
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1517_
timestamp 1667941163
transform 1 0 2024 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1517__85
timestamp 1667941163
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1518__86
timestamp 1667941163
transform 1 0 47748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1518_
timestamp 1667941163
transform 1 0 46460 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1519__87
timestamp 1667941163
transform 1 0 47472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1519_
timestamp 1667941163
transform 1 0 46460 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1520__88
timestamp 1667941163
transform 1 0 47748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1520_
timestamp 1667941163
transform 1 0 46460 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1521__89
timestamp 1667941163
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1521_
timestamp 1667941163
transform 1 0 2116 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1522_
timestamp 1667941163
transform 1 0 13616 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1522__90
timestamp 1667941163
transform 1 0 12880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1523__91
timestamp 1667941163
transform 1 0 44712 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1523_
timestamp 1667941163
transform 1 0 42780 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1524__92
timestamp 1667941163
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1524_
timestamp 1667941163
transform 1 0 12972 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1525__93
timestamp 1667941163
transform 1 0 35604 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1525_
timestamp 1667941163
transform 1 0 35512 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1526__94
timestamp 1667941163
transform 1 0 14352 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1526_
timestamp 1667941163
transform 1 0 14260 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1527_
timestamp 1667941163
transform 1 0 46460 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1527__95
timestamp 1667941163
transform 1 0 47748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1667941163
transform 1 0 2208 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1528__96
timestamp 1667941163
transform 1 0 2208 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1529__97
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1530__98
timestamp 1667941163
transform 1 0 23828 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1667941163
transform 1 0 24564 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1531__99
timestamp 1667941163
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1667941163
transform 1 0 24748 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1667941163
transform 1 0 45356 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1532__100
timestamp 1667941163
transform 1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1533__101
timestamp 1667941163
transform 1 0 47012 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1667941163
transform 1 0 46460 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1534__102
timestamp 1667941163
transform 1 0 28888 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1667941163
transform 1 0 29440 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1535__103
timestamp 1667941163
transform 1 0 41584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1667941163
transform 1 0 42596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1536__104
timestamp 1667941163
transform 1 0 47748 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1667941163
transform 1 0 46460 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1537__105
timestamp 1667941163
transform 1 0 7176 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1667941163
transform 1 0 1840 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1538__106
timestamp 1667941163
transform 1 0 40940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1667941163
transform 1 0 40480 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1539__107
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1540__108
timestamp 1667941163
transform 1 0 45816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1667941163
transform 1 0 45356 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1541__109
timestamp 1667941163
transform 1 0 10488 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1667941163
transform 1 0 10396 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1542__110
timestamp 1667941163
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1543__111
timestamp 1667941163
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1667941163
transform 1 0 2024 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1544__112
timestamp 1667941163
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1667941163
transform 1 0 2024 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36064 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1667941163
transform 1 0 28612 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1667941163
transform 1 0 31188 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1667941163
transform 1 0 26036 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1667941163
transform 1 0 31188 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1667941163
transform 1 0 36432 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1667941163
transform 1 0 41584 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1667941163
transform 1 0 39008 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1667941163
transform 1 0 41584 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 27784 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 7820 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 48116 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 48116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 9108 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1667941163
transform 1 0 47472 0 1 7616
box -38 -48 958 592
<< labels >>
flabel metal3 s 200 46188 800 46428 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 15446 200 15558 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 27682 49200 27794 49800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s -10 49200 102 49800 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 49200 42108 49800 42348 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 23818 200 23930 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 18666 49200 18778 49800 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 49200 44148 49800 44388 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 49200 4028 49800 4268 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 10294 49200 10406 49800 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 12226 49200 12338 49800 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 43138 200 43250 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 200 16268 800 16508 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 200 29188 800 29428 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 200 18988 800 19228 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 49200 15588 49800 15828 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 9006 49200 9118 49800 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 6430 49200 6542 49800 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 37342 200 37454 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 36698 200 36810 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 49200 10828 49800 11068 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 32834 200 32946 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 49578 49200 49690 49800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 16090 200 16202 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 49200 19668 49800 19908 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 200 44148 800 44388 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 30902 200 31014 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 200 25788 800 26028 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 37986 49200 38098 49800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 43138 49200 43250 49800 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 49200 31228 49800 31468 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 44426 49200 44538 49800 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 28970 49200 29082 49800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 49200 30548 49800 30788 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 49200 48228 49800 48468 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 200 30548 800 30788 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 200 21028 800 21268 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 49200 33268 49800 33508 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 8362 49200 8474 49800 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 26394 200 26506 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal bidirectional
flabel metal3 s 200 16948 800 17188 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal bidirectional
flabel metal3 s 49200 28508 49800 28748 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal bidirectional
flabel metal3 s 49200 14908 49800 15148 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal bidirectional
flabel metal3 s 49200 13548 49800 13788 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal bidirectional
flabel metal3 s 200 4708 800 4948 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal bidirectional
flabel metal2 s 14158 49200 14270 49800 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal bidirectional
flabel metal3 s 49200 1988 49800 2228 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal bidirectional
flabel metal2 s 13514 200 13626 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal bidirectional
flabel metal2 s 36054 49200 36166 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal bidirectional
flabel metal2 s 14802 49200 14914 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal bidirectional
flabel metal2 s 39274 200 39386 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal bidirectional
flabel metal3 s 49200 21708 49800 21948 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal bidirectional
flabel metal2 s 1922 49200 2034 49800 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal bidirectional
flabel metal2 s 5142 200 5254 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal bidirectional
flabel metal2 s 25106 49200 25218 49800 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal bidirectional
flabel metal2 s 25750 49200 25862 49800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal bidirectional
flabel metal2 s 47646 200 47758 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal bidirectional
flabel metal3 s 49200 39388 49800 39628 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal bidirectional
flabel metal2 s 29614 49200 29726 49800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal bidirectional
flabel metal2 s 41850 200 41962 800 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal bidirectional
flabel metal3 s 49200 32588 49800 32828 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal bidirectional
flabel metal2 s 41850 49200 41962 49800 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal bidirectional
flabel metal2 s 2566 49200 2678 49800 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal bidirectional
flabel metal2 s 41206 200 41318 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal bidirectional
flabel metal3 s 200 25108 800 25348 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal bidirectional
flabel metal2 s 48934 200 49046 800 0 FreeSans 448 90 0 0 io_oeb[33]
port 65 nsew signal bidirectional
flabel metal2 s 10938 49200 11050 49800 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal bidirectional
flabel metal3 s 200 21708 800 21948 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal bidirectional
flabel metal3 s 200 11508 800 11748 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal bidirectional
flabel metal3 s 200 18308 800 18548 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal bidirectional
flabel metal2 s 25750 200 25862 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal bidirectional
flabel metal3 s 49200 -52 49800 188 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal bidirectional
flabel metal3 s 200 32588 800 32828 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal bidirectional
flabel metal3 s 49200 17628 49800 17868 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal bidirectional
flabel metal2 s 12870 49200 12982 49800 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal bidirectional
flabel metal2 s 4498 200 4610 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal bidirectional
flabel metal2 s 10938 200 11050 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal bidirectional
flabel metal3 s 49200 46868 49800 47108 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal bidirectional
flabel metal3 s 49200 27828 49800 28068 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal bidirectional
flabel metal3 s 200 2668 800 2908 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal bidirectional
flabel metal3 s 200 7428 800 7668 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal bidirectional
flabel metal2 s 40562 200 40674 800 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal bidirectional
flabel metal3 s 49200 40068 49800 40308 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal bidirectional
flabel metal3 s 200 41428 800 41668 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal bidirectional
flabel metal3 s 49200 26468 49800 26708 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal bidirectional
flabel metal2 s 46358 49200 46470 49800 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal bidirectional
flabel metal2 s 47002 200 47114 800 0 FreeSans 448 90 0 0 io_out[18]
port 86 nsew signal bidirectional
flabel metal3 s 200 23748 800 23988 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal bidirectional
flabel metal2 s 33478 49200 33590 49800 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal bidirectional
flabel metal2 s 40562 49200 40674 49800 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal bidirectional
flabel metal3 s 200 40748 800 40988 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal bidirectional
flabel metal2 s 32190 200 32302 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal bidirectional
flabel metal3 s 49200 22388 49800 22628 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal bidirectional
flabel metal2 s 27682 200 27794 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal bidirectional
flabel metal2 s 36698 49200 36810 49800 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal bidirectional
flabel metal3 s 200 5388 800 5628 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal bidirectional
flabel metal2 s 38630 49200 38742 49800 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal bidirectional
flabel metal2 s 17378 200 17490 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal bidirectional
flabel metal3 s 49200 1308 49800 1548 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal bidirectional
flabel metal2 s 7074 200 7186 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal bidirectional
flabel metal3 s 200 6748 800 6988 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal bidirectional
flabel metal3 s 200 14228 800 14468 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal bidirectional
flabel metal3 s 200 47548 800 47788 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal bidirectional
flabel metal3 s 49200 6748 49800 6988 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal bidirectional
flabel metal3 s 49200 41428 49800 41668 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal bidirectional
flabel metal3 s 49200 38028 49800 38268 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal bidirectional
flabel metal2 s 15446 49200 15558 49800 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal bidirectional
flabel metal3 s 49200 44828 49800 45068 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal bidirectional
flabel metal3 s 200 43468 800 43708 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal bidirectional
flabel metal3 s 49200 29188 49800 29428 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal bidirectional
flabel metal2 s 23174 49200 23286 49800 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal bidirectional
flabel metal2 s 48290 49200 48402 49800 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal bidirectional
flabel metal3 s 200 20348 800 20588 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal bidirectional
flabel metal2 s 19310 200 19422 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal bidirectional
flabel metal3 s 200 14908 800 15148 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal bidirectional
flabel metal3 s 49200 8108 49800 8348 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 21886 200 21998 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 49200 6068 49800 6308 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 200 37348 800 37588 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 34122 200 34234 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 200 13548 800 13788 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 16734 49200 16846 49800 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 31546 49200 31658 49800 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 23818 49200 23930 49800 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal2 s 43782 200 43894 800 0 FreeSans 448 90 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 17378 49200 17490 49800 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 19954 200 20066 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 200 36668 800 36908 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 48934 49200 49046 49800 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 49200 8788 49800 9028 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 200 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 14158 200 14270 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 200 38708 800 38948 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 49200 3348 49800 3588 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 28970 200 29082 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 200 33948 800 34188 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal2 s 1278 49200 1390 49800 0 FreeSans 448 90 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 11582 200 11694 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 200 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal2 s 38630 200 38742 800 0 FreeSans 448 90 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 200 31908 800 32148 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 42494 49200 42606 49800 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 49200 24428 49800 24668 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 19310 49200 19422 49800 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 200 23068 800 23308 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 20598 49200 20710 49800 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 200 34628 800 34868 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 7718 200 7830 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal bidirectional
flabel metal3 s 49200 12188 49800 12428 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal bidirectional
flabel metal2 s 22530 200 22642 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal bidirectional
flabel metal3 s 49200 46188 49800 46428 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal bidirectional
flabel metal2 s 4498 49200 4610 49800 0 FreeSans 448 90 0 0 la1_data_out[13]
port 151 nsew signal bidirectional
flabel metal2 s 27038 49200 27150 49800 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal bidirectional
flabel metal3 s 200 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal bidirectional
flabel metal3 s 49200 16948 49800 17188 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal bidirectional
flabel metal3 s 49200 35988 49800 36228 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal bidirectional
flabel metal2 s 5786 49200 5898 49800 0 FreeSans 448 90 0 0 la1_data_out[18]
port 156 nsew signal bidirectional
flabel metal3 s 49200 25788 49800 26028 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal bidirectional
flabel metal3 s 200 45508 800 45748 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal bidirectional
flabel metal3 s 200 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal bidirectional
flabel metal3 s 49200 42788 49800 43028 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal bidirectional
flabel metal2 s 30258 49200 30370 49800 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal bidirectional
flabel metal2 s 12870 200 12982 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal bidirectional
flabel metal3 s 49200 18988 49800 19228 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal bidirectional
flabel metal3 s 200 3348 800 3588 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal bidirectional
flabel metal3 s 49200 5388 49800 5628 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal bidirectional
flabel metal3 s 200 48228 800 48468 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal bidirectional
flabel metal2 s 45070 200 45182 800 0 FreeSans 448 90 0 0 la1_data_out[28]
port 167 nsew signal bidirectional
flabel metal2 s 6430 200 6542 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal bidirectional
flabel metal2 s 20598 200 20710 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal bidirectional
flabel metal3 s 49200 12868 49800 13108 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal bidirectional
flabel metal3 s 49200 48908 49800 49148 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal bidirectional
flabel metal3 s 200 9468 800 9708 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal bidirectional
flabel metal2 s 45714 200 45826 800 0 FreeSans 448 90 0 0 la1_data_out[4]
port 173 nsew signal bidirectional
flabel metal2 s 3210 200 3322 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal bidirectional
flabel metal3 s 49200 20348 49800 20588 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal bidirectional
flabel metal2 s 634 200 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal bidirectional
flabel metal3 s 49200 37348 49800 37588 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal bidirectional
flabel metal2 s 47002 49200 47114 49800 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal bidirectional
flabel metal2 s 49578 200 49690 800 0 FreeSans 448 90 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 45070 49200 45182 49800 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 200 27828 800 28068 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 200 29868 800 30108 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 30258 200 30370 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 200 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 35410 200 35522 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 200 35988 800 36228 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal2 s 3854 49200 3966 49800 0 FreeSans 448 90 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 21886 49200 21998 49800 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 200 27148 800 27388 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 9006 200 9118 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 2566 200 2678 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 32190 49200 32302 49800 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 21242 49200 21354 49800 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 24462 200 24574 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 39918 49200 40030 49800 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 49200 10148 49800 10388 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 200 39388 800 39628 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 49200 35308 49800 35548 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 9650 200 9762 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 18022 200 18134 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 200 8108 800 8348 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 49200 34628 49800 34868 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 28326 200 28438 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 35410 49200 35522 49800 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 34122 49200 34234 49800 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 200 49588 800 49828 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal2 s 7718 49200 7830 49800 0 FreeSans 448 90 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 34766 200 34878 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 200 12188 800 12428 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 200 42788 800 43028 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 49200 23748 49800 23988 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
rlabel metal1 24978 47328 24978 47328 0 vccd1
rlabel metal1 24978 46784 24978 46784 0 vssd1
rlabel metal2 33810 23970 33810 23970 0 _0000_
rlabel metal1 34495 24786 34495 24786 0 _0001_
rlabel metal1 33994 22202 33994 22202 0 _0002_
rlabel metal1 37991 21930 37991 21930 0 _0003_
rlabel metal1 38732 24378 38732 24378 0 _0004_
rlabel metal1 40613 22610 40613 22610 0 _0005_
rlabel via1 42913 24786 42913 24786 0 _0006_
rlabel metal1 42810 24106 42810 24106 0 _0007_
rlabel metal2 31878 20706 31878 20706 0 _0008_
rlabel metal1 29808 20570 29808 20570 0 _0009_
rlabel metal1 31310 23018 31310 23018 0 _0010_
rlabel metal1 33074 28186 33074 28186 0 _0011_
rlabel metal1 30176 27098 30176 27098 0 _0012_
rlabel metal2 29854 25058 29854 25058 0 _0013_
rlabel metal2 30406 23970 30406 23970 0 _0014_
rlabel metal1 29746 21930 29746 21930 0 _0015_
rlabel metal2 38042 28662 38042 28662 0 _0016_
rlabel metal1 39785 25874 39785 25874 0 _0017_
rlabel metal2 39146 27846 39146 27846 0 _0018_
rlabel metal2 42366 28254 42366 28254 0 _0019_
rlabel via1 43557 25874 43557 25874 0 _0020_
rlabel metal2 43194 27846 43194 27846 0 _0021_
rlabel metal1 46271 27030 46271 27030 0 _0022_
rlabel metal1 45632 28730 45632 28730 0 _0023_
rlabel metal1 33488 32402 33488 32402 0 _0024_
rlabel metal2 33534 26758 33534 26758 0 _0025_
rlabel metal2 36202 26486 36202 26486 0 _0026_
rlabel metal2 32890 20230 32890 20230 0 _0027_
rlabel metal2 35374 20706 35374 20706 0 _0028_
rlabel metal1 37950 20026 37950 20026 0 _0029_
rlabel metal2 41354 20230 41354 20230 0 _0030_
rlabel metal2 43010 20706 43010 20706 0 _0031_
rlabel metal2 42090 21760 42090 21760 0 _0032_
rlabel via1 24881 32810 24881 32810 0 _0033_
rlabel metal1 35553 30634 35553 30634 0 _0034_
rlabel metal1 29803 29138 29803 29138 0 _0035_
rlabel metal2 27186 29410 27186 29410 0 _0036_
rlabel metal2 23414 30022 23414 30022 0 _0037_
rlabel via1 24881 27438 24881 27438 0 _0038_
rlabel metal2 23414 25670 23414 25670 0 _0039_
rlabel via1 24973 23086 24973 23086 0 _0040_
rlabel metal1 24600 21522 24600 21522 0 _0041_
rlabel metal2 27554 20536 27554 20536 0 _0042_
rlabel metal1 37664 37842 37664 37842 0 _0043_
rlabel metal2 27186 33762 27186 33762 0 _0044_
rlabel metal1 37352 32266 37352 32266 0 _0045_
rlabel metal2 37490 33762 37490 33762 0 _0046_
rlabel metal1 37945 30702 37945 30702 0 _0047_
rlabel metal1 41768 32538 41768 32538 0 _0048_
rlabel metal1 43086 30294 43086 30294 0 _0049_
rlabel metal1 46920 31178 46920 31178 0 _0050_
rlabel metal2 42918 35462 42918 35462 0 _0051_
rlabel metal1 47140 35054 47140 35054 0 _0052_
rlabel metal1 25944 31450 25944 31450 0 _0053_
rlabel metal1 29194 31382 29194 31382 0 _0054_
rlabel via1 31597 29614 31597 29614 0 _0055_
rlabel metal2 33166 30498 33166 30498 0 _0056_
rlabel metal1 29389 32470 29389 32470 0 _0057_
rlabel metal2 28934 34374 28934 34374 0 _0058_
rlabel metal1 29164 35258 29164 35258 0 _0059_
rlabel metal1 31045 34578 31045 34578 0 _0060_
rlabel metal1 40015 37910 40015 37910 0 _0061_
rlabel metal1 32384 32538 32384 32538 0 _0062_
rlabel metal1 39049 39406 39049 39406 0 _0063_
rlabel metal1 35829 36074 35829 36074 0 _0064_
rlabel via1 34541 33558 34541 33558 0 _0065_
rlabel metal2 35742 34374 35742 34374 0 _0066_
rlabel metal1 32568 35258 32568 35258 0 _0067_
rlabel metal1 31947 37094 31947 37094 0 _0068_
rlabel via1 31137 38318 31137 38318 0 _0069_
rlabel metal1 33207 37910 33207 37910 0 _0070_
rlabel metal1 34771 36822 34771 36822 0 _0071_
rlabel metal1 23996 42262 23996 42262 0 _0072_
rlabel metal1 27871 36754 27871 36754 0 _0073_
rlabel metal1 24318 35734 24318 35734 0 _0074_
rlabel metal1 24140 34578 24140 34578 0 _0075_
rlabel via1 23869 37910 23869 37910 0 _0076_
rlabel metal1 23920 39610 23920 39610 0 _0077_
rlabel metal1 24196 40698 24196 40698 0 _0078_
rlabel metal2 26450 39202 26450 39202 0 _0079_
rlabel viali 25893 35054 25893 35054 0 _0080_
rlabel metal1 27360 42194 27360 42194 0 _0081_
rlabel metal1 28469 38998 28469 38998 0 _0082_
rlabel metal1 28458 40086 28458 40086 0 _0083_
rlabel metal1 27181 41514 27181 41514 0 _0084_
rlabel metal2 29026 42670 29026 42670 0 _0085_
rlabel metal1 30171 42670 30171 42670 0 _0086_
rlabel metal1 32936 42330 32936 42330 0 _0087_
rlabel metal1 32103 41514 32103 41514 0 _0088_
rlabel via1 28377 37842 28377 37842 0 _0089_
rlabel metal1 24134 41514 24134 41514 0 _0090_
rlabel metal1 33667 40018 33667 40018 0 _0091_
rlabel metal1 33529 40494 33529 40494 0 _0092_
rlabel metal1 34541 42194 34541 42194 0 _0093_
rlabel metal2 35926 42874 35926 42874 0 _0094_
rlabel metal1 36703 41514 36703 41514 0 _0095_
rlabel metal1 38394 41174 38394 41174 0 _0096_
rlabel metal1 39095 40086 39095 40086 0 _0097_
rlabel via1 35737 38998 35737 38998 0 _0098_
rlabel metal2 42642 37026 42642 37026 0 _0099_
rlabel metal1 43546 37910 43546 37910 0 _0100_
rlabel metal1 45662 38998 45662 38998 0 _0101_
rlabel metal1 45126 39610 45126 39610 0 _0102_
rlabel metal1 45075 41174 45075 41174 0 _0103_
rlabel metal1 43516 41786 43516 41786 0 _0104_
rlabel via1 41165 40494 41165 40494 0 _0105_
rlabel metal1 42688 39610 42688 39610 0 _0106_
rlabel metal1 41763 38250 41763 38250 0 _0107_
rlabel metal1 5014 44812 5014 44812 0 _0108_
rlabel metal1 3634 17646 3634 17646 0 _0109_
rlabel metal2 20746 3774 20746 3774 0 _0110_
rlabel metal1 4416 2414 4416 2414 0 _0111_
rlabel metal1 2530 4080 2530 4080 0 _0112_
rlabel metal1 2852 19822 2852 19822 0 _0113_
rlabel metal1 40710 3094 40710 3094 0 _0114_
rlabel metal1 2530 21386 2530 21386 0 _0115_
rlabel metal1 5796 44778 5796 44778 0 _0116_
rlabel metal1 2714 16626 2714 16626 0 _0117_
rlabel metal1 5658 2414 5658 2414 0 _0118_
rlabel metal1 2898 21522 2898 21522 0 _0119_
rlabel metal1 44022 21998 44022 21998 0 _0120_
rlabel metal2 44114 23460 44114 23460 0 _0121_
rlabel metal1 41032 18258 41032 18258 0 _0122_
rlabel metal1 37766 18768 37766 18768 0 _0123_
rlabel metal2 36570 19482 36570 19482 0 _0124_
rlabel metal2 36846 18972 36846 18972 0 _0125_
rlabel metal1 36846 22746 36846 22746 0 _0126_
rlabel metal1 36984 24174 36984 24174 0 _0127_
rlabel metal1 38364 23834 38364 23834 0 _0128_
rlabel metal1 37076 23018 37076 23018 0 _0129_
rlabel metal1 36616 24174 36616 24174 0 _0130_
rlabel metal2 36938 23562 36938 23562 0 _0131_
rlabel metal2 36662 23290 36662 23290 0 _0132_
rlabel metal1 37858 23120 37858 23120 0 _0133_
rlabel metal1 37858 22746 37858 22746 0 _0134_
rlabel metal2 37398 22814 37398 22814 0 _0135_
rlabel metal1 39882 22746 39882 22746 0 _0136_
rlabel metal2 43838 23290 43838 23290 0 _0137_
rlabel metal2 44482 22780 44482 22780 0 _0138_
rlabel metal2 38364 31756 38364 31756 0 _0139_
rlabel metal2 34362 21216 34362 21216 0 _0140_
rlabel metal1 26450 20910 26450 20910 0 _0141_
rlabel via1 27646 22627 27646 22627 0 _0142_
rlabel metal1 24288 23834 24288 23834 0 _0143_
rlabel metal1 24334 25466 24334 25466 0 _0144_
rlabel metal2 26634 27268 26634 27268 0 _0145_
rlabel metal1 27600 27302 27600 27302 0 _0146_
rlabel metal2 27462 26554 27462 26554 0 _0147_
rlabel metal2 28198 26044 28198 26044 0 _0148_
rlabel metal2 28566 26010 28566 26010 0 _0149_
rlabel metal1 28336 24378 28336 24378 0 _0150_
rlabel metal1 27968 23290 27968 23290 0 _0151_
rlabel metal2 27646 24956 27646 24956 0 _0152_
rlabel metal2 28106 25942 28106 25942 0 _0153_
rlabel metal1 26956 26350 26956 26350 0 _0154_
rlabel metal1 27186 25908 27186 25908 0 _0155_
rlabel metal1 27186 24208 27186 24208 0 _0156_
rlabel metal1 27324 23086 27324 23086 0 _0157_
rlabel metal1 27232 22746 27232 22746 0 _0158_
rlabel metal2 32522 24038 32522 24038 0 _0159_
rlabel metal1 32200 38930 32200 38930 0 _0160_
rlabel metal2 33534 33694 33534 33694 0 _0161_
rlabel metal1 42964 41582 42964 41582 0 _0162_
rlabel metal1 45954 37366 45954 37366 0 _0163_
rlabel metal1 45726 30702 45726 30702 0 _0164_
rlabel metal2 45218 29988 45218 29988 0 _0165_
rlabel metal1 44068 28730 44068 28730 0 _0166_
rlabel metal1 43746 29648 43746 29648 0 _0167_
rlabel metal2 41998 29750 41998 29750 0 _0168_
rlabel metal2 43286 29376 43286 29376 0 _0169_
rlabel metal1 40664 29818 40664 29818 0 _0170_
rlabel metal2 40250 29920 40250 29920 0 _0171_
rlabel metal2 40066 30192 40066 30192 0 _0172_
rlabel metal1 37628 32402 37628 32402 0 _0173_
rlabel metal1 39422 29818 39422 29818 0 _0174_
rlabel metal1 39146 30260 39146 30260 0 _0175_
rlabel metal1 40480 30362 40480 30362 0 _0176_
rlabel metal2 41170 30498 41170 30498 0 _0177_
rlabel metal2 42366 29920 42366 29920 0 _0178_
rlabel metal1 43102 29172 43102 29172 0 _0179_
rlabel metal1 43010 29274 43010 29274 0 _0180_
rlabel metal2 45586 30396 45586 30396 0 _0181_
rlabel metal1 45783 37094 45783 37094 0 _0182_
rlabel metal1 46092 37434 46092 37434 0 _0183_
rlabel metal2 35466 24582 35466 24582 0 _0184_
rlabel metal1 34546 22134 34546 22134 0 _0185_
rlabel metal1 34454 22066 34454 22066 0 _0186_
rlabel metal1 38180 21658 38180 21658 0 _0187_
rlabel metal2 41170 26656 41170 26656 0 _0188_
rlabel metal2 38318 23290 38318 23290 0 _0189_
rlabel metal2 38870 24786 38870 24786 0 _0190_
rlabel metal1 40480 23222 40480 23222 0 _0191_
rlabel metal1 41170 24582 41170 24582 0 _0192_
rlabel metal2 41998 24480 41998 24480 0 _0193_
rlabel metal2 42182 25092 42182 25092 0 _0194_
rlabel metal2 42274 24786 42274 24786 0 _0195_
rlabel metal2 29946 20876 29946 20876 0 _0196_
rlabel metal1 30958 22474 30958 22474 0 _0197_
rlabel metal2 31970 27642 31970 27642 0 _0198_
rlabel metal1 32430 27574 32430 27574 0 _0199_
rlabel metal1 32844 28050 32844 28050 0 _0200_
rlabel metal1 30360 26962 30360 26962 0 _0201_
rlabel metal1 30038 26996 30038 26996 0 _0202_
rlabel metal1 31050 24922 31050 24922 0 _0203_
rlabel metal1 30452 24786 30452 24786 0 _0204_
rlabel metal2 30498 23868 30498 23868 0 _0205_
rlabel metal2 31234 24378 31234 24378 0 _0206_
rlabel metal1 29670 22542 29670 22542 0 _0207_
rlabel metal1 40250 26384 40250 26384 0 _0208_
rlabel metal2 39238 28118 39238 28118 0 _0209_
rlabel metal1 41768 27438 41768 27438 0 _0210_
rlabel metal1 42274 27642 42274 27642 0 _0211_
rlabel metal1 42044 28526 42044 28526 0 _0212_
rlabel metal1 43654 26384 43654 26384 0 _0213_
rlabel metal2 43378 27132 43378 27132 0 _0214_
rlabel metal1 45954 27472 45954 27472 0 _0215_
rlabel metal2 45954 28288 45954 28288 0 _0216_
rlabel metal1 46644 27642 46644 27642 0 _0217_
rlabel via1 45773 28186 45773 28186 0 _0218_
rlabel metal2 34178 33082 34178 33082 0 _0219_
rlabel metal1 36708 28526 36708 28526 0 _0220_
rlabel metal1 35374 28594 35374 28594 0 _0221_
rlabel metal1 35558 28628 35558 28628 0 _0222_
rlabel metal2 35374 29580 35374 29580 0 _0223_
rlabel metal1 40756 21998 40756 21998 0 _0224_
rlabel metal1 35006 20468 35006 20468 0 _0225_
rlabel metal1 33718 26384 33718 26384 0 _0226_
rlabel metal1 35650 29104 35650 29104 0 _0227_
rlabel metal1 35604 18802 35604 18802 0 _0228_
rlabel metal1 35972 19822 35972 19822 0 _0229_
rlabel metal2 36386 25670 36386 25670 0 _0230_
rlabel metal1 35098 27472 35098 27472 0 _0231_
rlabel metal1 35558 26010 35558 26010 0 _0232_
rlabel metal1 37352 25874 37352 25874 0 _0233_
rlabel metal1 36662 25908 36662 25908 0 _0234_
rlabel metal1 38134 33456 38134 33456 0 _0235_
rlabel metal2 35374 28169 35374 28169 0 _0236_
rlabel metal1 36064 19414 36064 19414 0 _0237_
rlabel metal2 35190 19380 35190 19380 0 _0238_
rlabel metal1 34454 19346 34454 19346 0 _0239_
rlabel metal1 33902 19278 33902 19278 0 _0240_
rlabel metal1 33764 19482 33764 19482 0 _0241_
rlabel metal1 34316 18938 34316 18938 0 _0242_
rlabel viali 35114 19346 35114 19346 0 _0243_
rlabel metal1 34592 20026 34592 20026 0 _0244_
rlabel metal1 35374 20026 35374 20026 0 _0245_
rlabel metal1 34914 20332 34914 20332 0 _0246_
rlabel metal3 33718 20604 33718 20604 0 _0247_
rlabel metal1 35604 19346 35604 19346 0 _0248_
rlabel metal2 38778 19074 38778 19074 0 _0249_
rlabel metal1 38640 18734 38640 18734 0 _0250_
rlabel metal2 38962 19142 38962 19142 0 _0251_
rlabel metal1 38732 19278 38732 19278 0 _0252_
rlabel metal1 38456 19482 38456 19482 0 _0253_
rlabel metal2 40250 18564 40250 18564 0 _0254_
rlabel metal1 39928 18802 39928 18802 0 _0255_
rlabel metal2 40618 19312 40618 19312 0 _0256_
rlabel metal2 41262 19652 41262 19652 0 _0257_
rlabel metal2 44022 19482 44022 19482 0 _0258_
rlabel metal2 44390 19074 44390 19074 0 _0259_
rlabel metal1 43608 19346 43608 19346 0 _0260_
rlabel metal1 40342 19346 40342 19346 0 _0261_
rlabel metal1 40158 19448 40158 19448 0 _0262_
rlabel metal2 43194 19652 43194 19652 0 _0263_
rlabel metal1 43378 20026 43378 20026 0 _0264_
rlabel metal1 44252 19278 44252 19278 0 _0265_
rlabel metal1 44252 21862 44252 21862 0 _0266_
rlabel metal1 41630 21624 41630 21624 0 _0267_
rlabel metal1 41860 21522 41860 21522 0 _0268_
rlabel metal1 39330 42126 39330 42126 0 _0269_
rlabel metal1 24426 33524 24426 33524 0 _0270_
rlabel metal1 35604 31790 35604 31790 0 _0271_
rlabel metal2 26634 30974 26634 30974 0 _0272_
rlabel metal1 27554 31314 27554 31314 0 _0273_
rlabel metal1 25898 32198 25898 32198 0 _0274_
rlabel metal1 26634 31824 26634 31824 0 _0275_
rlabel metal1 27232 21522 27232 21522 0 _0276_
rlabel metal1 29670 28968 29670 28968 0 _0277_
rlabel metal2 30774 28934 30774 28934 0 _0278_
rlabel metal1 26726 32198 26726 32198 0 _0279_
rlabel metal1 26266 31926 26266 31926 0 _0280_
rlabel metal1 23184 20434 23184 20434 0 _0281_
rlabel metal1 26358 28730 26358 28730 0 _0282_
rlabel metal1 26358 29580 26358 29580 0 _0283_
rlabel metal2 26818 28764 26818 28764 0 _0284_
rlabel metal1 27508 28526 27508 28526 0 _0285_
rlabel metal2 27646 28934 27646 28934 0 _0286_
rlabel metal2 26634 30090 26634 30090 0 _0287_
rlabel metal2 24610 29308 24610 29308 0 _0288_
rlabel metal1 24656 28458 24656 28458 0 _0289_
rlabel metal1 24334 28730 24334 28730 0 _0290_
rlabel metal2 24518 28458 24518 28458 0 _0291_
rlabel metal2 23966 29376 23966 29376 0 _0292_
rlabel metal2 23414 27744 23414 27744 0 _0293_
rlabel metal1 25362 28118 25362 28118 0 _0294_
rlabel metal2 23874 27999 23874 27999 0 _0295_
rlabel metal2 22678 27914 22678 27914 0 _0296_
rlabel metal1 22908 27574 22908 27574 0 _0297_
rlabel metal2 23782 27710 23782 27710 0 _0298_
rlabel metal1 23046 25262 23046 25262 0 _0299_
rlabel metal2 22402 24242 22402 24242 0 _0300_
rlabel metal1 23184 24786 23184 24786 0 _0301_
rlabel metal1 23506 24684 23506 24684 0 _0302_
rlabel metal1 23782 24922 23782 24922 0 _0303_
rlabel metal1 23000 23630 23000 23630 0 _0304_
rlabel metal1 23644 23154 23644 23154 0 _0305_
rlabel metal1 24196 23290 24196 23290 0 _0306_
rlabel metal2 25530 23868 25530 23868 0 _0307_
rlabel metal1 23368 22610 23368 22610 0 _0308_
rlabel metal1 23092 21998 23092 21998 0 _0309_
rlabel metal1 23460 21862 23460 21862 0 _0310_
rlabel metal1 24104 23698 24104 23698 0 _0311_
rlabel metal1 23598 21964 23598 21964 0 _0312_
rlabel metal1 24058 20910 24058 20910 0 _0313_
rlabel metal2 23782 21318 23782 21318 0 _0314_
rlabel metal2 26266 21250 26266 21250 0 _0315_
rlabel metal2 26358 20570 26358 20570 0 _0316_
rlabel metal1 26634 20536 26634 20536 0 _0317_
rlabel metal2 27462 20876 27462 20876 0 _0318_
rlabel metal2 36938 38012 36938 38012 0 _0319_
rlabel metal2 27370 33932 27370 33932 0 _0320_
rlabel metal1 39882 35700 39882 35700 0 _0321_
rlabel metal2 39606 35836 39606 35836 0 _0322_
rlabel metal2 39698 36074 39698 36074 0 _0323_
rlabel metal2 40710 35836 40710 35836 0 _0324_
rlabel metal2 38594 35258 38594 35258 0 _0325_
rlabel metal1 39146 32980 39146 32980 0 _0326_
rlabel metal2 38042 34680 38042 34680 0 _0327_
rlabel metal1 37904 31994 37904 31994 0 _0328_
rlabel metal2 40986 36380 40986 36380 0 _0329_
rlabel metal1 40296 32946 40296 32946 0 _0330_
rlabel metal1 40848 34374 40848 34374 0 _0331_
rlabel metal1 40250 34000 40250 34000 0 _0332_
rlabel metal1 39514 34612 39514 34612 0 _0333_
rlabel metal1 38456 33490 38456 33490 0 _0334_
rlabel metal2 38962 34238 38962 34238 0 _0335_
rlabel metal1 38916 33626 38916 33626 0 _0336_
rlabel metal1 37950 33524 37950 33524 0 _0337_
rlabel metal1 40158 34578 40158 34578 0 _0338_
rlabel metal1 39468 31790 39468 31790 0 _0339_
rlabel metal2 40066 32028 40066 32028 0 _0340_
rlabel metal1 40388 31994 40388 31994 0 _0341_
rlabel metal1 40986 31790 40986 31790 0 _0342_
rlabel metal1 38824 32742 38824 32742 0 _0343_
rlabel metal2 41262 33014 41262 33014 0 _0344_
rlabel metal1 41032 32946 41032 32946 0 _0345_
rlabel metal2 41170 32844 41170 32844 0 _0346_
rlabel metal2 40894 32164 40894 32164 0 _0347_
rlabel metal1 40618 31450 40618 31450 0 _0348_
rlabel metal1 42550 31722 42550 31722 0 _0349_
rlabel metal1 44114 32946 44114 32946 0 _0350_
rlabel metal1 44068 31994 44068 31994 0 _0351_
rlabel metal2 44850 32640 44850 32640 0 _0352_
rlabel metal1 43424 32198 43424 32198 0 _0353_
rlabel metal1 45356 32946 45356 32946 0 _0354_
rlabel metal1 45770 32334 45770 32334 0 _0355_
rlabel metal1 46828 31314 46828 31314 0 _0356_
rlabel metal1 47150 31416 47150 31416 0 _0357_
rlabel metal2 44022 35122 44022 35122 0 _0358_
rlabel metal1 44666 35802 44666 35802 0 _0359_
rlabel metal2 44206 35530 44206 35530 0 _0360_
rlabel metal1 45448 31994 45448 31994 0 _0361_
rlabel metal2 44574 33830 44574 33830 0 _0362_
rlabel metal1 43286 35156 43286 35156 0 _0363_
rlabel metal1 43516 34714 43516 34714 0 _0364_
rlabel metal1 45862 34612 45862 34612 0 _0365_
rlabel metal2 45954 34816 45954 34816 0 _0366_
rlabel metal1 46736 34442 46736 34442 0 _0367_
rlabel metal1 46920 34714 46920 34714 0 _0368_
rlabel metal1 24748 31314 24748 31314 0 _0369_
rlabel metal1 33350 35020 33350 35020 0 _0370_
rlabel metal2 30130 31110 30130 31110 0 _0371_
rlabel metal2 31694 30396 31694 30396 0 _0372_
rlabel metal1 33028 30226 33028 30226 0 _0373_
rlabel metal2 30590 32436 30590 32436 0 _0374_
rlabel metal1 29118 34000 29118 34000 0 _0375_
rlabel metal1 29210 35088 29210 35088 0 _0376_
rlabel metal1 31280 35054 31280 35054 0 _0377_
rlabel metal1 39744 38318 39744 38318 0 _0378_
rlabel metal2 32522 33184 32522 33184 0 _0379_
rlabel metal1 32476 32402 32476 32402 0 _0380_
rlabel metal2 31786 32130 31786 32130 0 _0381_
rlabel metal1 31372 32878 31372 32878 0 _0382_
rlabel via1 32811 32470 32811 32470 0 _0383_
rlabel metal2 40250 41548 40250 41548 0 _0384_
rlabel metal1 36984 35666 36984 35666 0 _0385_
rlabel metal2 34362 34170 34362 34170 0 _0386_
rlabel metal1 35604 33966 35604 33966 0 _0387_
rlabel metal1 32706 35088 32706 35088 0 _0388_
rlabel metal2 32890 38522 32890 38522 0 _0389_
rlabel metal1 32062 36890 32062 36890 0 _0390_
rlabel metal1 31326 37978 31326 37978 0 _0391_
rlabel metal1 33396 38318 33396 38318 0 _0392_
rlabel via1 34738 35802 34738 35802 0 _0393_
rlabel metal2 34914 36023 34914 36023 0 _0394_
rlabel metal2 36478 36924 36478 36924 0 _0395_
rlabel metal1 35926 36618 35926 36618 0 _0396_
rlabel metal2 36202 37026 36202 37026 0 _0397_
rlabel metal2 23690 42908 23690 42908 0 _0398_
rlabel metal2 28474 36618 28474 36618 0 _0399_
rlabel metal2 23414 36618 23414 36618 0 _0400_
rlabel metal2 24058 36346 24058 36346 0 _0401_
rlabel metal1 24426 37434 24426 37434 0 _0402_
rlabel metal1 24058 39440 24058 39440 0 _0403_
rlabel metal1 24058 40528 24058 40528 0 _0404_
rlabel metal2 26634 39372 26634 39372 0 _0405_
rlabel metal1 25589 36890 25589 36890 0 _0406_
rlabel metal1 25668 36754 25668 36754 0 _0407_
rlabel metal2 27554 36550 27554 36550 0 _0408_
rlabel metal2 26266 37774 26266 37774 0 _0409_
rlabel via1 26279 36822 26279 36822 0 _0410_
rlabel metal2 27370 43452 27370 43452 0 _0411_
rlabel metal1 28290 38318 28290 38318 0 _0412_
rlabel metal1 30084 39610 30084 39610 0 _0413_
rlabel metal2 37674 41888 37674 41888 0 _0414_
rlabel metal2 28934 42194 28934 42194 0 _0415_
rlabel metal2 29210 42364 29210 42364 0 _0416_
rlabel metal1 30314 42262 30314 42262 0 _0417_
rlabel metal1 33166 42160 33166 42160 0 _0418_
rlabel metal1 32614 41242 32614 41242 0 _0419_
rlabel metal1 30514 40426 30514 40426 0 _0420_
rlabel metal1 28474 39440 28474 39440 0 _0421_
rlabel metal1 30314 39950 30314 39950 0 _0422_
rlabel metal2 30866 40460 30866 40460 0 _0423_
rlabel metal1 29647 39338 29647 39338 0 _0424_
rlabel metal2 23598 42636 23598 42636 0 _0425_
rlabel metal1 32706 39406 32706 39406 0 _0426_
rlabel metal1 34132 39610 34132 39610 0 _0427_
rlabel metal1 35328 41786 35328 41786 0 _0428_
rlabel metal2 36110 42806 36110 42806 0 _0429_
rlabel metal1 36938 42228 36938 42228 0 _0430_
rlabel metal2 38594 41990 38594 41990 0 _0431_
rlabel metal1 39422 40460 39422 40460 0 _0432_
rlabel metal1 36213 40426 36213 40426 0 _0433_
rlabel viali 35374 40040 35374 40040 0 _0434_
rlabel metal2 35466 39746 35466 39746 0 _0435_
rlabel metal2 36662 40460 36662 40460 0 _0436_
rlabel metal1 35995 40086 35995 40086 0 _0437_
rlabel metal1 42366 35802 42366 35802 0 _0438_
rlabel metal2 44298 37536 44298 37536 0 _0439_
rlabel metal2 45586 38726 45586 38726 0 _0440_
rlabel metal2 45402 39610 45402 39610 0 _0441_
rlabel metal1 45494 41582 45494 41582 0 _0442_
rlabel metal1 43424 41582 43424 41582 0 _0443_
rlabel metal2 41814 40562 41814 40562 0 _0444_
rlabel metal2 42550 40154 42550 40154 0 _0445_
rlabel metal2 42826 39066 42826 39066 0 _0446_
rlabel metal1 42734 38250 42734 38250 0 _0447_
rlabel metal1 43562 39032 43562 39032 0 _0448_
rlabel metal1 43332 38998 43332 38998 0 _0449_
rlabel metal1 43401 38250 43401 38250 0 _0450_
rlabel metal1 8096 3094 8096 3094 0 _0451_
rlabel metal2 2438 44574 2438 44574 0 _0452_
rlabel metal1 20332 3094 20332 3094 0 _0453_
rlabel metal2 2346 8670 2346 8670 0 _0454_
rlabel metal2 45402 3468 45402 3468 0 _0455_
rlabel metal2 4002 3978 4002 3978 0 _0456_
rlabel metal2 46690 20060 46690 20060 0 _0457_
rlabel metal1 3358 2346 3358 2346 0 _0458_
rlabel metal1 47288 37162 47288 37162 0 _0459_
rlabel metal1 45908 45050 45908 45050 0 _0460_
rlabel metal2 46690 11356 46690 11356 0 _0461_
rlabel metal2 22218 3230 22218 3230 0 _0462_
rlabel metal1 46736 45526 46736 45526 0 _0463_
rlabel metal1 4554 45050 4554 45050 0 _0464_
rlabel metal2 27002 46308 27002 46308 0 _0465_
rlabel metal1 2070 2924 2070 2924 0 _0466_
rlabel metal2 47886 16354 47886 16354 0 _0467_
rlabel metal1 47288 36210 47288 36210 0 _0468_
rlabel metal2 6670 45730 6670 45730 0 _0469_
rlabel metal2 47150 25296 47150 25296 0 _0470_
rlabel metal2 2898 9758 2898 9758 0 _0471_
rlabel metal1 47288 42738 47288 42738 0 _0472_
rlabel metal1 29900 45594 29900 45594 0 _0473_
rlabel metal1 12282 2482 12282 2482 0 _0474_
rlabel metal1 46920 18802 46920 18802 0 _0475_
rlabel metal1 2208 4250 2208 4250 0 _0476_
rlabel metal2 46690 5916 46690 5916 0 _0477_
rlabel metal2 1794 46444 1794 46444 0 _0478_
rlabel metal2 45126 3502 45126 3502 0 _0479_
rlabel metal1 6026 3434 6026 3434 0 _0480_
rlabel metal1 46920 12274 46920 12274 0 _0481_
rlabel metal2 45586 46546 45586 46546 0 _0482_
rlabel metal2 47150 43554 47150 43554 0 _0483_
rlabel metal2 33258 46308 33258 46308 0 _0484_
rlabel metal1 7038 3910 7038 3910 0 _0485_
rlabel metal2 2622 43554 2622 43554 0 _0486_
rlabel metal1 47288 29546 47288 29546 0 _0487_
rlabel metal2 22954 46308 22954 46308 0 _0488_
rlabel metal1 48116 46138 48116 46138 0 _0489_
rlabel metal2 2530 20196 2530 20196 0 _0490_
rlabel metal1 19550 2482 19550 2482 0 _0491_
rlabel metal2 2254 15198 2254 15198 0 _0492_
rlabel metal1 47288 26418 47288 26418 0 _0493_
rlabel metal1 1794 3604 1794 3604 0 _0494_
rlabel metal1 2277 7922 2277 7922 0 _0495_
rlabel metal2 40250 2652 40250 2652 0 _0496_
rlabel metal2 46874 38114 46874 38114 0 _0497_
rlabel metal2 28474 23188 28474 23188 0 _0498_
rlabel metal1 45678 23290 45678 23290 0 _0499_
rlabel metal1 46046 24378 46046 24378 0 _0500_
rlabel metal2 45862 3944 45862 3944 0 _0501_
rlabel metal1 2392 23290 2392 23290 0 _0502_
rlabel metal2 40342 45458 40342 45458 0 _0503_
rlabel metal2 2438 40868 2438 40868 0 _0504_
rlabel metal2 32522 3230 32522 3230 0 _0505_
rlabel metal2 47150 22882 47150 22882 0 _0506_
rlabel metal2 27646 2788 27646 2788 0 _0507_
rlabel metal1 37168 45526 37168 45526 0 _0508_
rlabel metal2 2898 6052 2898 6052 0 _0509_
rlabel metal1 39008 46138 39008 46138 0 _0510_
rlabel metal2 17066 3230 17066 3230 0 _0511_
rlabel metal2 38594 3230 38594 3230 0 _0512_
rlabel metal2 4094 7140 4094 7140 0 _0513_
rlabel metal1 2346 14042 2346 14042 0 _0514_
rlabel metal2 6762 46750 6762 46750 0 _0515_
rlabel metal2 47886 6562 47886 6562 0 _0516_
rlabel metal1 47288 41650 47288 41650 0 _0517_
rlabel metal1 47288 39474 47288 39474 0 _0518_
rlabel metal1 15686 46070 15686 46070 0 _0519_
rlabel metal1 46598 44506 46598 44506 0 _0520_
rlabel metal1 25714 3434 25714 3434 0 _0521_
rlabel metal2 39422 3808 39422 3808 0 _0522_
rlabel metal1 42228 45526 42228 45526 0 _0523_
rlabel metal2 24978 3230 24978 3230 0 _0524_
rlabel metal1 46598 4522 46598 4522 0 _0525_
rlabel metal2 2438 32674 2438 32674 0 _0526_
rlabel metal1 47288 17714 47288 17714 0 _0527_
rlabel metal2 12466 46002 12466 46002 0 _0528_
rlabel metal2 4922 4828 4922 4828 0 _0529_
rlabel metal2 10534 3740 10534 3740 0 _0530_
rlabel metal1 2576 17238 2576 17238 0 _0531_
rlabel metal2 47886 28322 47886 28322 0 _0532_
rlabel metal2 46690 14620 46690 14620 0 _0533_
rlabel metal1 46920 13362 46920 13362 0 _0534_
rlabel metal2 4094 5406 4094 5406 0 _0535_
rlabel metal1 13478 45526 13478 45526 0 _0536_
rlabel metal2 43010 3196 43010 3196 0 _0537_
rlabel metal2 13202 3502 13202 3502 0 _0538_
rlabel metal2 35742 45730 35742 45730 0 _0539_
rlabel metal1 14076 45866 14076 45866 0 _0540_
rlabel metal2 47150 21794 47150 21794 0 _0541_
rlabel metal1 2116 44506 2116 44506 0 _0542_
rlabel metal1 5014 3094 5014 3094 0 _0543_
rlabel metal1 24656 45594 24656 45594 0 _0544_
rlabel metal1 25162 45594 25162 45594 0 _0545_
rlabel metal1 47426 2618 47426 2618 0 _0546_
rlabel metal1 47288 40562 47288 40562 0 _0547_
rlabel metal1 29394 46138 29394 46138 0 _0548_
rlabel metal2 42826 3230 42826 3230 0 _0549_
rlabel metal2 47886 32674 47886 32674 0 _0550_
rlabel metal1 3082 46614 3082 46614 0 _0551_
rlabel metal2 41446 3264 41446 3264 0 _0552_
rlabel metal1 2116 24922 2116 24922 0 _0553_
rlabel metal2 44574 4964 44574 4964 0 _0554_
rlabel metal2 10626 45730 10626 45730 0 _0555_
rlabel metal1 2346 21658 2346 21658 0 _0556_
rlabel metal2 2346 11492 2346 11492 0 _0557_
rlabel metal1 2484 17850 2484 17850 0 _0558_
rlabel metal1 2346 42670 2346 42670 0 active
rlabel metal1 37904 36822 37904 36822 0 clknet_0_wb_clk_i
rlabel metal1 26910 21012 26910 21012 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 32338 20672 32338 20672 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 26082 33184 26082 33184 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 33902 42398 33902 42398 0 clknet_3_3__leaf_wb_clk_i
rlabel metal1 37306 32844 37306 32844 0 clknet_3_4__leaf_wb_clk_i
rlabel metal1 40526 20468 40526 20468 0 clknet_3_5__leaf_wb_clk_i
rlabel metal1 36938 41582 36938 41582 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 46966 33456 46966 33456 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 28014 48161 28014 48161 0 io_in[10]
rlabel metal2 46 49038 46 49038 0 io_in[11]
rlabel metal2 48346 43299 48346 43299 0 io_in[12]
rlabel metal2 23874 1588 23874 1588 0 io_in[13]
rlabel metal2 48346 33677 48346 33677 0 io_in[8]
rlabel metal1 8878 47022 8878 47022 0 io_in[9]
rlabel metal2 26450 2166 26450 2166 0 io_oeb[0]
rlabel metal3 1740 17068 1740 17068 0 io_oeb[10]
rlabel metal3 48814 28628 48814 28628 0 io_oeb[11]
rlabel metal3 48814 15028 48814 15028 0 io_oeb[12]
rlabel metal3 48814 13668 48814 13668 0 io_oeb[13]
rlabel metal2 2806 4981 2806 4981 0 io_oeb[14]
rlabel metal2 14214 47338 14214 47338 0 io_oeb[15]
rlabel metal1 44666 2312 44666 2312 0 io_oeb[16]
rlabel metal2 13570 1860 13570 1860 0 io_oeb[17]
rlabel metal2 36110 47644 36110 47644 0 io_oeb[18]
rlabel metal2 14858 47644 14858 47644 0 io_oeb[19]
rlabel metal2 39330 2370 39330 2370 0 io_oeb[1]
rlabel metal3 48860 21828 48860 21828 0 io_oeb[20]
rlabel metal1 2484 46410 2484 46410 0 io_oeb[21]
rlabel metal2 5198 1860 5198 1860 0 io_oeb[22]
rlabel metal2 25162 47644 25162 47644 0 io_oeb[23]
rlabel metal2 25806 47882 25806 47882 0 io_oeb[24]
rlabel metal2 47702 2404 47702 2404 0 io_oeb[25]
rlabel metal3 48814 39508 48814 39508 0 io_oeb[26]
rlabel metal1 29854 46478 29854 46478 0 io_oeb[27]
rlabel metal2 41906 1860 41906 1860 0 io_oeb[28]
rlabel metal3 48860 32708 48860 32708 0 io_oeb[29]
rlabel metal1 43102 46444 43102 46444 0 io_oeb[2]
rlabel metal1 2714 46478 2714 46478 0 io_oeb[30]
rlabel metal2 41262 2166 41262 2166 0 io_oeb[31]
rlabel metal3 1740 25228 1740 25228 0 io_oeb[32]
rlabel metal2 48990 2948 48990 2948 0 io_oeb[33]
rlabel metal1 11040 46002 11040 46002 0 io_oeb[34]
rlabel metal3 1740 21828 1740 21828 0 io_oeb[35]
rlabel via2 2806 11645 2806 11645 0 io_oeb[36]
rlabel metal2 2806 18309 2806 18309 0 io_oeb[37]
rlabel metal2 25806 1860 25806 1860 0 io_oeb[3]
rlabel metal3 48860 68 48860 68 0 io_oeb[4]
rlabel metal3 1740 32708 1740 32708 0 io_oeb[5]
rlabel metal3 48814 17748 48814 17748 0 io_oeb[6]
rlabel metal2 12926 47882 12926 47882 0 io_oeb[7]
rlabel metal2 4554 1571 4554 1571 0 io_oeb[8]
rlabel metal2 10994 2166 10994 2166 0 io_oeb[9]
rlabel metal3 48768 46988 48768 46988 0 io_out[0]
rlabel metal3 48814 27948 48814 27948 0 io_out[10]
rlabel metal2 2806 3179 2806 3179 0 io_out[11]
rlabel metal2 2990 7735 2990 7735 0 io_out[12]
rlabel metal2 40618 1622 40618 1622 0 io_out[13]
rlabel metal3 48722 40188 48722 40188 0 io_out[14]
rlabel metal3 2108 41548 2108 41548 0 io_out[15]
rlabel metal3 48722 26588 48722 26588 0 io_out[16]
rlabel metal2 45816 45540 45816 45540 0 io_out[17]
rlabel metal2 47058 2098 47058 2098 0 io_out[18]
rlabel metal2 2806 23749 2806 23749 0 io_out[19]
rlabel metal2 33534 47882 33534 47882 0 io_out[1]
rlabel metal2 40618 47644 40618 47644 0 io_out[20]
rlabel metal3 1740 40868 1740 40868 0 io_out[21]
rlabel metal2 32246 1860 32246 1860 0 io_out[22]
rlabel metal3 48860 22508 48860 22508 0 io_out[23]
rlabel metal2 27738 1860 27738 1860 0 io_out[24]
rlabel metal1 37950 46444 37950 46444 0 io_out[25]
rlabel metal2 2990 5865 2990 5865 0 io_out[26]
rlabel metal1 40250 46444 40250 46444 0 io_out[27]
rlabel metal2 17434 1860 17434 1860 0 io_out[28]
rlabel metal1 40250 2924 40250 2924 0 io_out[29]
rlabel metal2 7130 1027 7130 1027 0 io_out[2]
rlabel metal2 2806 7089 2806 7089 0 io_out[30]
rlabel metal3 1740 14348 1740 14348 0 io_out[31]
rlabel metal3 2108 47668 2108 47668 0 io_out[32]
rlabel metal3 48814 6868 48814 6868 0 io_out[33]
rlabel metal3 48814 41548 48814 41548 0 io_out[34]
rlabel metal3 48768 38148 48768 38148 0 io_out[35]
rlabel metal2 15502 47882 15502 47882 0 io_out[36]
rlabel metal3 48814 44948 48814 44948 0 io_out[37]
rlabel metal3 1740 43588 1740 43588 0 io_out[3]
rlabel metal3 48860 29308 48860 29308 0 io_out[4]
rlabel metal2 23230 47882 23230 47882 0 io_out[5]
rlabel metal2 48346 47950 48346 47950 0 io_out[6]
rlabel metal3 1740 20468 1740 20468 0 io_out[7]
rlabel metal2 19366 1027 19366 1027 0 io_out[8]
rlabel metal3 1740 15028 1740 15028 0 io_out[9]
rlabel metal2 47518 8075 47518 8075 0 la1_data_in[0]
rlabel metal2 7774 1761 7774 1761 0 la1_data_out[0]
rlabel metal3 48124 12308 48124 12308 0 la1_data_out[10]
rlabel metal2 22586 1860 22586 1860 0 la1_data_out[11]
rlabel metal3 48124 46308 48124 46308 0 la1_data_out[12]
rlabel metal2 4738 47889 4738 47889 0 la1_data_out[13]
rlabel metal1 27646 46444 27646 46444 0 la1_data_out[14]
rlabel metal3 1786 1428 1786 1428 0 la1_data_out[15]
rlabel metal3 48814 17068 48814 17068 0 la1_data_out[16]
rlabel metal3 48814 36108 48814 36108 0 la1_data_out[17]
rlabel metal2 5842 47644 5842 47644 0 la1_data_out[18]
rlabel metal3 48308 25908 48308 25908 0 la1_data_out[19]
rlabel metal3 1740 45628 1740 45628 0 la1_data_out[1]
rlabel metal2 2990 9877 2990 9877 0 la1_data_out[20]
rlabel metal3 48814 42908 48814 42908 0 la1_data_out[21]
rlabel metal1 30360 46002 30360 46002 0 la1_data_out[22]
rlabel metal2 12926 1622 12926 1622 0 la1_data_out[23]
rlabel metal3 48814 19108 48814 19108 0 la1_data_out[24]
rlabel metal2 2990 4063 2990 4063 0 la1_data_out[25]
rlabel metal3 48814 5508 48814 5508 0 la1_data_out[26]
rlabel metal2 2806 47175 2806 47175 0 la1_data_out[27]
rlabel metal2 45126 1860 45126 1860 0 la1_data_out[28]
rlabel metal1 6578 3570 6578 3570 0 la1_data_out[29]
rlabel metal2 20654 1860 20654 1860 0 la1_data_out[2]
rlabel metal3 48814 12988 48814 12988 0 la1_data_out[30]
rlabel metal3 48308 49028 48308 49028 0 la1_data_out[31]
rlabel metal2 2806 8993 2806 8993 0 la1_data_out[3]
rlabel metal2 45770 1622 45770 1622 0 la1_data_out[4]
rlabel metal2 3266 1792 3266 1792 0 la1_data_out[5]
rlabel metal3 48814 20468 48814 20468 0 la1_data_out[6]
rlabel metal2 690 1622 690 1622 0 la1_data_out[7]
rlabel metal3 48814 37468 48814 37468 0 la1_data_out[8]
rlabel metal2 47058 47678 47058 47678 0 la1_data_out[9]
rlabel metal1 2162 42534 2162 42534 0 net1
rlabel metal2 2254 44812 2254 44812 0 net10
rlabel metal1 45402 4012 45402 4012 0 net100
rlabel metal2 46506 40732 46506 40732 0 net101
rlabel metal1 29302 46546 29302 46546 0 net102
rlabel metal2 42642 3468 42642 3468 0 net103
rlabel metal1 47242 32946 47242 32946 0 net104
rlabel metal1 1886 46614 1886 46614 0 net105
rlabel metal2 40526 3740 40526 3740 0 net106
rlabel metal2 1610 25500 1610 25500 0 net107
rlabel metal1 45402 5236 45402 5236 0 net108
rlabel metal2 10442 46172 10442 46172 0 net109
rlabel metal1 19964 2958 19964 2958 0 net11
rlabel metal1 1978 21522 1978 21522 0 net110
rlabel metal1 2070 11764 2070 11764 0 net111
rlabel metal2 2070 18496 2070 18496 0 net112
rlabel metal2 2162 8704 2162 8704 0 net12
rlabel metal1 44850 2482 44850 2482 0 net13
rlabel metal1 4002 2618 4002 2618 0 net14
rlabel metal1 46506 19924 46506 19924 0 net15
rlabel metal1 1610 2346 1610 2346 0 net16
rlabel metal1 46506 37162 46506 37162 0 net17
rlabel metal2 45770 46172 45770 46172 0 net18
rlabel metal1 46506 11220 46506 11220 0 net19
rlabel metal1 27508 43758 27508 43758 0 net2
rlabel metal2 22034 3264 22034 3264 0 net20
rlabel metal1 45172 45390 45172 45390 0 net21
rlabel metal2 4186 46784 4186 46784 0 net22
rlabel metal2 27186 46784 27186 46784 0 net23
rlabel metal1 1886 3060 1886 3060 0 net24
rlabel metal2 46506 16796 46506 16796 0 net25
rlabel metal2 46506 36380 46506 36380 0 net26
rlabel metal1 5612 46002 5612 46002 0 net27
rlabel metal1 47426 24718 47426 24718 0 net28
rlabel metal2 2162 9792 2162 9792 0 net29
rlabel metal2 7866 45118 7866 45118 0 net3
rlabel metal1 46276 42670 46276 42670 0 net30
rlabel metal1 29854 46002 29854 46002 0 net31
rlabel metal1 11914 2516 11914 2516 0 net32
rlabel metal1 46506 18836 46506 18836 0 net33
rlabel metal1 1840 4114 1840 4114 0 net34
rlabel metal2 47978 5406 47978 5406 0 net35
rlabel metal1 2346 45866 2346 45866 0 net36
rlabel metal2 44942 3264 44942 3264 0 net37
rlabel metal1 6210 3638 6210 3638 0 net38
rlabel metal1 46506 12308 46506 12308 0 net39
rlabel metal1 40066 42228 40066 42228 0 net4
rlabel metal1 44712 46070 44712 46070 0 net40
rlabel metal1 46874 43826 46874 43826 0 net41
rlabel metal1 32982 46580 32982 46580 0 net42
rlabel metal1 6946 2482 6946 2482 0 net43
rlabel metal1 1840 43282 1840 43282 0 net44
rlabel metal1 46874 29682 46874 29682 0 net45
rlabel metal2 22494 46784 22494 46784 0 net46
rlabel metal1 45034 46546 45034 46546 0 net47
rlabel metal2 2070 20672 2070 20672 0 net48
rlabel metal1 19412 2414 19412 2414 0 net49
rlabel metal1 24610 2482 24610 2482 0 net5
rlabel metal1 2024 14994 2024 14994 0 net50
rlabel metal2 47978 26078 47978 26078 0 net51
rlabel metal1 1656 3570 1656 3570 0 net52
rlabel metal1 1978 6970 1978 6970 0 net53
rlabel metal2 40066 3536 40066 3536 0 net54
rlabel metal1 46920 3570 46920 3570 0 net55
rlabel metal2 2070 23936 2070 23936 0 net56
rlabel metal1 40296 45458 40296 45458 0 net57
rlabel metal2 2070 41344 2070 41344 0 net58
rlabel metal1 32108 3026 32108 3026 0 net59
rlabel metal2 48162 34850 48162 34850 0 net6
rlabel metal1 47978 22644 47978 22644 0 net60
rlabel metal2 27462 3264 27462 3264 0 net61
rlabel metal1 37030 46478 37030 46478 0 net62
rlabel metal1 2254 5882 2254 5882 0 net63
rlabel metal2 39790 46784 39790 46784 0 net64
rlabel metal2 16882 3264 16882 3264 0 net65
rlabel metal2 38410 3264 38410 3264 0 net66
rlabel metal1 2070 7276 2070 7276 0 net67
rlabel metal1 1978 13906 1978 13906 0 net68
rlabel metal2 6578 46784 6578 46784 0 net69
rlabel metal2 9154 45084 9154 45084 0 net7
rlabel metal1 46690 6834 46690 6834 0 net70
rlabel metal2 46506 41820 46506 41820 0 net71
rlabel metal2 46506 39644 46506 39644 0 net72
rlabel metal1 14490 46580 14490 46580 0 net73
rlabel metal2 46506 45084 46506 45084 0 net74
rlabel metal2 25898 3740 25898 3740 0 net75
rlabel metal1 38824 2618 38824 2618 0 net76
rlabel metal2 42642 46784 42642 46784 0 net77
rlabel metal2 24794 3468 24794 3468 0 net78
rlabel metal2 47978 4386 47978 4386 0 net79
rlabel metal1 46920 7854 46920 7854 0 net8
rlabel metal1 1978 32946 1978 32946 0 net80
rlabel metal1 47242 17170 47242 17170 0 net81
rlabel metal1 12190 46580 12190 46580 0 net82
rlabel metal1 4508 4590 4508 4590 0 net83
rlabel metal1 10442 3026 10442 3026 0 net84
rlabel metal1 2208 16762 2208 16762 0 net85
rlabel metal1 47242 28594 47242 28594 0 net86
rlabel metal1 46506 14484 46506 14484 0 net87
rlabel metal1 46506 13396 46506 13396 0 net88
rlabel metal1 2162 5270 2162 5270 0 net89
rlabel metal2 7590 3468 7590 3468 0 net9
rlabel metal1 13524 45458 13524 45458 0 net90
rlabel metal1 42826 2516 42826 2516 0 net91
rlabel metal2 13018 3264 13018 3264 0 net92
rlabel metal2 35558 46172 35558 46172 0 net93
rlabel metal1 14444 46002 14444 46002 0 net94
rlabel metal1 47978 21556 47978 21556 0 net95
rlabel metal1 2392 42738 2392 42738 0 net96
rlabel metal2 4186 3264 4186 3264 0 net97
rlabel metal1 24334 45934 24334 45934 0 net98
rlabel metal1 24794 46580 24794 46580 0 net99
rlabel metal2 44298 38522 44298 38522 0 rgb_mixer.debounce0_a.button_hist\[0\]
rlabel metal1 45172 38318 45172 38318 0 rgb_mixer.debounce0_a.button_hist\[1\]
rlabel metal1 44206 38862 44206 38862 0 rgb_mixer.debounce0_a.button_hist\[2\]
rlabel metal2 45310 40324 45310 40324 0 rgb_mixer.debounce0_a.button_hist\[3\]
rlabel metal1 42734 41616 42734 41616 0 rgb_mixer.debounce0_a.button_hist\[4\]
rlabel metal1 43562 41106 43562 41106 0 rgb_mixer.debounce0_a.button_hist\[5\]
rlabel metal1 42780 41106 42780 41106 0 rgb_mixer.debounce0_a.button_hist\[6\]
rlabel metal2 42918 40256 42918 40256 0 rgb_mixer.debounce0_a.button_hist\[7\]
rlabel metal1 40262 37162 40262 37162 0 rgb_mixer.debounce0_a.debounced
rlabel metal1 27002 41786 27002 41786 0 rgb_mixer.debounce0_b.button_hist\[0\]
rlabel metal2 34546 40290 34546 40290 0 rgb_mixer.debounce0_b.button_hist\[1\]
rlabel metal1 34868 41582 34868 41582 0 rgb_mixer.debounce0_b.button_hist\[2\]
rlabel metal1 35420 41990 35420 41990 0 rgb_mixer.debounce0_b.button_hist\[3\]
rlabel metal1 37352 42126 37352 42126 0 rgb_mixer.debounce0_b.button_hist\[4\]
rlabel metal1 37996 41446 37996 41446 0 rgb_mixer.debounce0_b.button_hist\[5\]
rlabel metal1 37352 40426 37352 40426 0 rgb_mixer.debounce0_b.button_hist\[6\]
rlabel metal2 37214 40256 37214 40256 0 rgb_mixer.debounce0_b.button_hist\[7\]
rlabel metal1 36800 39066 36800 39066 0 rgb_mixer.debounce0_b.debounced
rlabel metal1 28428 40698 28428 40698 0 rgb_mixer.debounce1_a.button_hist\[0\]
rlabel metal1 29762 40460 29762 40460 0 rgb_mixer.debounce1_a.button_hist\[1\]
rlabel metal1 29992 40154 29992 40154 0 rgb_mixer.debounce1_a.button_hist\[2\]
rlabel metal1 28566 40528 28566 40528 0 rgb_mixer.debounce1_a.button_hist\[3\]
rlabel metal2 29854 42636 29854 42636 0 rgb_mixer.debounce1_a.button_hist\[4\]
rlabel metal1 31004 41106 31004 41106 0 rgb_mixer.debounce1_a.button_hist\[5\]
rlabel metal1 32706 42534 32706 42534 0 rgb_mixer.debounce1_a.button_hist\[6\]
rlabel metal1 30774 41514 30774 41514 0 rgb_mixer.debounce1_a.button_hist\[7\]
rlabel metal1 30222 37978 30222 37978 0 rgb_mixer.debounce1_a.debounced
rlabel metal1 27692 35462 27692 35462 0 rgb_mixer.debounce1_b.button_hist\[0\]
rlabel metal2 27370 36108 27370 36108 0 rgb_mixer.debounce1_b.button_hist\[1\]
rlabel metal2 26082 36873 26082 36873 0 rgb_mixer.debounce1_b.button_hist\[2\]
rlabel metal2 26174 37077 26174 37077 0 rgb_mixer.debounce1_b.button_hist\[3\]
rlabel metal2 25622 39134 25622 39134 0 rgb_mixer.debounce1_b.button_hist\[4\]
rlabel metal2 25070 40290 25070 40290 0 rgb_mixer.debounce1_b.button_hist\[5\]
rlabel metal2 25622 40460 25622 40460 0 rgb_mixer.debounce1_b.button_hist\[6\]
rlabel metal2 25714 39168 25714 39168 0 rgb_mixer.debounce1_b.button_hist\[7\]
rlabel metal1 26680 35258 26680 35258 0 rgb_mixer.debounce1_b.debounced
rlabel metal1 38042 36686 38042 36686 0 rgb_mixer.debounce2_a.button_hist\[0\]
rlabel metal1 34546 35700 34546 35700 0 rgb_mixer.debounce2_a.button_hist\[1\]
rlabel metal1 35052 35462 35052 35462 0 rgb_mixer.debounce2_a.button_hist\[2\]
rlabel metal1 34592 34714 34592 34714 0 rgb_mixer.debounce2_a.button_hist\[3\]
rlabel metal2 33442 36176 33442 36176 0 rgb_mixer.debounce2_a.button_hist\[4\]
rlabel metal1 33074 37400 33074 37400 0 rgb_mixer.debounce2_a.button_hist\[5\]
rlabel metal1 32706 38420 32706 38420 0 rgb_mixer.debounce2_a.button_hist\[6\]
rlabel metal1 33672 37230 33672 37230 0 rgb_mixer.debounce2_a.button_hist\[7\]
rlabel metal1 35742 36856 35742 36856 0 rgb_mixer.debounce2_a.debounced
rlabel metal2 29762 31212 29762 31212 0 rgb_mixer.debounce2_b.button_hist\[0\]
rlabel metal1 32062 31110 32062 31110 0 rgb_mixer.debounce2_b.button_hist\[1\]
rlabel metal1 32246 30226 32246 30226 0 rgb_mixer.debounce2_b.button_hist\[2\]
rlabel metal1 30774 31382 30774 31382 0 rgb_mixer.debounce2_b.button_hist\[3\]
rlabel metal2 29854 33252 29854 33252 0 rgb_mixer.debounce2_b.button_hist\[4\]
rlabel metal2 31142 33558 31142 33558 0 rgb_mixer.debounce2_b.button_hist\[5\]
rlabel metal2 30590 35292 30590 35292 0 rgb_mixer.debounce2_b.button_hist\[6\]
rlabel metal2 31786 34170 31786 34170 0 rgb_mixer.debounce2_b.button_hist\[7\]
rlabel metal1 33488 32742 33488 32742 0 rgb_mixer.debounce2_b.debounced
rlabel metal1 38686 31824 38686 31824 0 rgb_mixer.enc0\[0\]
rlabel metal1 40894 33932 40894 33932 0 rgb_mixer.enc0\[1\]
rlabel metal1 39100 32402 39100 32402 0 rgb_mixer.enc0\[2\]
rlabel metal2 41354 32521 41354 32521 0 rgb_mixer.enc0\[3\]
rlabel metal1 44390 32334 44390 32334 0 rgb_mixer.enc0\[4\]
rlabel metal2 45126 29852 45126 29852 0 rgb_mixer.enc0\[5\]
rlabel metal1 44804 33966 44804 33966 0 rgb_mixer.enc0\[6\]
rlabel metal1 46460 34578 46460 34578 0 rgb_mixer.enc0\[7\]
rlabel metal1 26726 28526 26726 28526 0 rgb_mixer.enc1\[0\]
rlabel metal2 27462 28288 27462 28288 0 rgb_mixer.enc1\[1\]
rlabel metal1 23828 26962 23828 26962 0 rgb_mixer.enc1\[2\]
rlabel metal1 25254 26928 25254 26928 0 rgb_mixer.enc1\[3\]
rlabel metal1 25024 25262 25024 25262 0 rgb_mixer.enc1\[4\]
rlabel metal1 25714 24208 25714 24208 0 rgb_mixer.enc1\[5\]
rlabel metal1 26128 21658 26128 21658 0 rgb_mixer.enc1\[6\]
rlabel metal2 28290 21318 28290 21318 0 rgb_mixer.enc1\[7\]
rlabel metal2 35374 25840 35374 25840 0 rgb_mixer.enc2\[0\]
rlabel metal1 35190 28628 35190 28628 0 rgb_mixer.enc2\[1\]
rlabel metal1 36478 19822 36478 19822 0 rgb_mixer.enc2\[2\]
rlabel metal1 36478 20400 36478 20400 0 rgb_mixer.enc2\[3\]
rlabel metal1 38962 19856 38962 19856 0 rgb_mixer.enc2\[4\]
rlabel metal2 41906 20026 41906 20026 0 rgb_mixer.enc2\[5\]
rlabel metal1 44896 21114 44896 21114 0 rgb_mixer.enc2\[6\]
rlabel metal1 39514 24038 39514 24038 0 rgb_mixer.enc2\[7\]
rlabel metal1 40756 37298 40756 37298 0 rgb_mixer.encoder0.old_a
rlabel metal2 40342 37434 40342 37434 0 rgb_mixer.encoder0.old_b
rlabel metal2 27094 32810 27094 32810 0 rgb_mixer.encoder1.old_a
rlabel metal1 26266 32300 26266 32300 0 rgb_mixer.encoder1.old_b
rlabel metal2 36202 30090 36202 30090 0 rgb_mixer.encoder2.old_a
rlabel metal1 35512 30226 35512 30226 0 rgb_mixer.encoder2.old_b
rlabel metal1 39652 29002 39652 29002 0 rgb_mixer.pwm0.count\[0\]
rlabel metal2 40250 28798 40250 28798 0 rgb_mixer.pwm0.count\[1\]
rlabel metal1 40066 28560 40066 28560 0 rgb_mixer.pwm0.count\[2\]
rlabel metal2 41538 28832 41538 28832 0 rgb_mixer.pwm0.count\[3\]
rlabel metal2 43930 28390 43930 28390 0 rgb_mixer.pwm0.count\[4\]
rlabel metal2 43746 27200 43746 27200 0 rgb_mixer.pwm0.count\[5\]
rlabel metal1 45724 27506 45724 27506 0 rgb_mixer.pwm0.count\[6\]
rlabel metal1 45954 28594 45954 28594 0 rgb_mixer.pwm0.count\[7\]
rlabel metal2 46138 38148 46138 38148 0 rgb_mixer.pwm0.out
rlabel metal1 31556 20434 31556 20434 0 rgb_mixer.pwm1.count\[0\]
rlabel metal1 31280 21114 31280 21114 0 rgb_mixer.pwm1.count\[1\]
rlabel metal1 30866 23766 30866 23766 0 rgb_mixer.pwm1.count\[2\]
rlabel metal2 32338 28220 32338 28220 0 rgb_mixer.pwm1.count\[3\]
rlabel metal2 27370 26044 27370 26044 0 rgb_mixer.pwm1.count\[4\]
rlabel metal2 27462 24922 27462 24922 0 rgb_mixer.pwm1.count\[5\]
rlabel via1 27648 24174 27648 24174 0 rgb_mixer.pwm1.count\[6\]
rlabel metal1 30590 22576 30590 22576 0 rgb_mixer.pwm1.count\[7\]
rlabel metal2 27738 23392 27738 23392 0 rgb_mixer.pwm1.out
rlabel metal1 34868 21930 34868 21930 0 rgb_mixer.pwm2.count\[0\]
rlabel metal1 35282 21998 35282 21998 0 rgb_mixer.pwm2.count\[1\]
rlabel metal1 34822 21998 34822 21998 0 rgb_mixer.pwm2.count\[2\]
rlabel metal1 37628 21454 37628 21454 0 rgb_mixer.pwm2.count\[3\]
rlabel metal2 39146 24650 39146 24650 0 rgb_mixer.pwm2.count\[4\]
rlabel metal1 39698 23018 39698 23018 0 rgb_mixer.pwm2.count\[5\]
rlabel metal1 41262 24752 41262 24752 0 rgb_mixer.pwm2.count\[6\]
rlabel metal1 38870 23664 38870 23664 0 rgb_mixer.pwm2.count\[7\]
rlabel metal2 45402 23154 45402 23154 0 rgb_mixer.pwm2.out
rlabel metal1 37766 24582 37766 24582 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
